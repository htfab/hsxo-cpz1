magic
tech sky130A
magscale 1 2
timestamp 1713788423
<< error_s >>
rect 1958 1573 1992 1956
rect 2080 1633 2138 1647
rect 2238 1633 2296 1647
rect 2154 1593 2222 1607
rect 2026 1579 2350 1593
rect 2138 1573 2260 1579
rect 2384 1573 2418 1956
rect 2568 1573 2602 1956
rect 2690 1633 2748 1647
rect 2848 1633 2906 1647
rect 2764 1593 2832 1607
rect 2636 1579 2960 1593
rect 2748 1573 2870 1579
rect 2994 1573 3028 1956
rect 3097 1573 3562 1682
rect 4841 1573 5304 1682
rect 5378 1573 5412 1956
rect 5500 1633 5558 1647
rect 5658 1633 5716 1647
rect 5574 1593 5642 1607
rect 5446 1579 5770 1593
rect 5558 1573 5680 1579
rect 5804 1573 5838 1956
rect 5988 1573 6022 1956
rect 6110 1633 6168 1647
rect 6268 1633 6326 1647
rect 6184 1593 6252 1607
rect 6056 1579 6380 1593
rect 6168 1573 6290 1579
rect 6414 1573 6448 1956
rect 797 1539 6823 1573
rect 1958 1510 1992 1539
rect 2138 1536 2238 1539
rect 2384 1510 2418 1539
rect 2568 1510 2602 1539
rect 2748 1536 2848 1539
rect 2994 1510 3028 1539
rect 3097 1474 3562 1539
rect 2982 1460 3562 1474
rect 3097 1446 3562 1460
rect 3010 1432 3562 1446
rect 3097 1286 3562 1432
rect 4841 1480 5304 1539
rect 5378 1510 5412 1539
rect 5558 1536 5658 1539
rect 5804 1510 5838 1539
rect 5988 1510 6022 1539
rect 6168 1536 6268 1539
rect 6414 1510 6448 1539
rect 4841 1474 5348 1480
rect 4841 1460 5428 1474
rect 4841 1452 5304 1460
rect 4841 1446 5320 1452
rect 4841 1432 5400 1446
rect 4841 1286 5304 1432
rect 2120 1282 2860 1286
rect 1910 930 3076 1282
rect 3080 930 5320 1286
rect 5540 1282 6290 1286
rect 6490 1282 6970 1286
rect 5241 886 5304 930
rect 5314 650 5320 930
rect 5241 566 5320 650
rect 5330 566 6970 1282
rect 5301 512 5314 566
rect 5300 112 5314 304
rect 6849 -2428 6883 0
rect 5874 -2462 7248 -2428
rect 6849 -2528 6883 -2462
rect 6832 -2539 6883 -2528
rect 6829 -2566 6883 -2539
rect 6884 -2566 6903 -2528
rect 6815 -2593 6883 -2566
rect 6895 -2593 6903 -2566
rect 6815 -2600 6903 -2593
rect 6906 -2600 6917 -2566
rect 6922 -2600 6941 -2566
rect 6829 -2625 6848 -2600
rect 6849 -2625 6903 -2600
rect 6826 -2659 6903 -2625
rect 6829 -3435 6917 -2659
rect 7114 -3244 7170 -3240
rect 7170 -3300 7226 -3284
rect 6829 -3447 6903 -3435
rect 6829 -3456 6848 -3447
rect 6849 -3456 6883 -3447
rect 6895 -3456 6903 -3447
rect 6829 -3494 6883 -3456
rect 6884 -3494 6903 -3456
rect 6815 -3528 6883 -3494
rect 6829 -3544 6848 -3528
rect 6829 -3555 6840 -3544
rect 6849 -3632 6883 -3528
rect 6895 -3555 6903 -3494
rect 6906 -3528 6917 -3494
rect 6922 -3528 6941 -3494
rect 5874 -3666 7248 -3632
rect 6849 -3754 6883 -3666
rect 6800 -5350 6970 -3754
rect 2030 -7244 2776 -7100
rect 1865 -7285 2776 -7244
rect 1865 -7302 3318 -7285
rect 2030 -7314 3318 -7302
rect 3420 -7314 5730 -7100
rect 2030 -7388 5730 -7314
rect 1890 -7608 5730 -7388
rect 2067 -7644 5730 -7608
rect 2067 -7654 2141 -7644
rect 2156 -7652 5730 -7644
rect 2156 -7654 4852 -7652
rect 1890 -7864 4852 -7654
rect 4858 -7750 4870 -7652
rect 1800 -7874 4852 -7864
rect 1800 -7944 2000 -7874
rect 1740 -7960 2000 -7944
rect 2030 -7910 4852 -7874
rect 2030 -7944 5017 -7910
rect 2030 -7960 3318 -7944
rect 1740 -7977 3318 -7960
rect 3441 -7968 5017 -7944
rect 1740 -8018 2776 -7977
rect 1740 -8024 2000 -8018
rect 1800 -8064 2000 -8024
rect 2030 -8274 2776 -8018
rect 2796 -8152 2830 -7977
rect 3441 -8133 4852 -7968
rect 5444 -7994 5730 -7652
rect 5806 -7910 5864 -7829
rect 5806 -7968 5895 -7910
rect 5641 -8133 5730 -7994
rect 0 -8800 70 -8798
rect 2190 -8800 2390 -8798
rect 0 -8944 70 -8804
rect 0 -9004 230 -8944
rect 30 -9144 230 -9004
<< dnwell >>
rect 760 -5240 6860 1550
rect 2110 -11280 5650 -7180
<< nwell >>
rect 650 930 6970 1660
rect 650 740 1570 930
rect 650 -2614 1370 740
rect 5314 196 6970 930
rect 5300 136 6970 196
rect 5530 130 6970 136
rect 650 -2814 1720 -2614
rect 650 -3160 1370 -2814
rect 650 -3360 4500 -3160
rect 650 -4920 966 -3360
rect 6654 -4920 6970 130
rect 650 -5020 970 -4920
rect 6650 -5020 6970 -4920
rect 650 -5350 6970 -5020
rect 2030 -7652 5730 -7100
rect 2030 -11074 2316 -7652
rect 5444 -11074 5730 -7652
rect 2030 -11360 5730 -11074
<< nsubdiff >>
rect 2067 -7157 5693 -7137
rect 2067 -7191 2147 -7157
rect 5613 -7191 5693 -7157
rect 2067 -7211 5693 -7191
rect 2067 -7217 2141 -7211
rect 2067 -11243 2087 -7217
rect 2121 -11243 2141 -7217
rect 2067 -11249 2141 -11243
rect 5619 -7217 5693 -7211
rect 5619 -11243 5639 -7217
rect 5673 -11243 5693 -7217
rect 5619 -11249 5693 -11243
rect 2067 -11269 5693 -11249
rect 2067 -11303 2147 -11269
rect 5613 -11303 5693 -11269
rect 2067 -11323 5693 -11303
<< mvnsubdiff >>
rect 717 1573 6903 1593
rect 717 1539 797 1573
rect 6823 1539 6903 1573
rect 717 1519 6903 1539
rect 717 1513 791 1519
rect 717 -5203 737 1513
rect 771 -5203 791 1513
rect 717 -5209 791 -5203
rect 6829 1513 6903 1519
rect 6829 -5203 6849 1513
rect 6883 -5203 6903 1513
rect 6829 -5209 6903 -5203
rect 717 -5229 6903 -5209
rect 717 -5263 797 -5229
rect 6823 -5263 6903 -5229
rect 717 -5283 6903 -5263
<< nsubdiffcont >>
rect 2147 -7191 5613 -7157
rect 2087 -11243 2121 -7217
rect 5639 -11243 5673 -7217
rect 2147 -11303 5613 -11269
<< mvnsubdiffcont >>
rect 797 1539 6823 1573
rect 737 -5203 771 1513
rect 6849 -5203 6883 1513
rect 797 -5263 6823 -5229
<< locali >>
rect 1076 5486 1264 5674
rect 737 1539 797 1573
rect 6823 1539 6883 1573
rect 737 1513 771 1539
rect 737 -5229 771 -5203
rect 6849 1513 6883 1539
rect 6849 -5229 6883 -5203
rect 737 -5263 797 -5229
rect 6823 -5263 6883 -5229
rect 2087 -7191 2147 -7157
rect 5613 -7191 5673 -7157
rect 2087 -7217 2121 -7191
rect 2087 -11269 2121 -11243
rect 5639 -7217 5673 -7191
rect 5639 -11269 5673 -11243
rect 2087 -11303 2147 -11269
rect 5613 -11303 5673 -11269
<< metal1 >>
rect 1070 5680 1270 5686
rect 1070 5474 1270 5480
rect -540 -544 -340 -538
rect -540 -8180 -340 -744
rect -140 -900 60 -898
rect -140 -904 70 -900
rect 60 -1104 70 -904
rect -140 -1110 70 -1104
rect -540 -8386 -340 -8380
rect -133 -8633 70 -1110
rect 284 -1474 290 -1274
rect 490 -1474 496 -1274
rect 290 -7698 490 -1474
rect 692 -1824 698 -1624
rect 898 -1824 904 -1624
rect -130 -8804 70 -8633
rect -136 -9004 -130 -8804
rect 70 -9004 76 -8804
rect 289 -10014 492 -7698
rect 284 -10214 290 -10014
rect 490 -10214 496 -10014
rect 290 -10744 490 -10738
rect 290 -11460 490 -10944
rect 698 -11098 898 -1824
rect 1050 -9314 1250 -9308
rect 698 -11104 900 -11098
rect 698 -11300 700 -11104
rect 700 -11310 900 -11304
rect 290 -11666 490 -11660
rect 1050 -11810 1250 -9514
rect 1044 -12010 1050 -11810
rect 1250 -12010 1256 -11810
<< via1 >>
rect 1070 5480 1270 5680
rect -540 -744 -340 -544
rect -140 -1104 60 -904
rect -540 -8380 -340 -8180
rect 290 -1474 490 -1274
rect 698 -1824 898 -1624
rect -130 -9004 70 -8804
rect 290 -10214 490 -10014
rect 290 -10944 490 -10744
rect 1050 -9514 1250 -9314
rect 700 -11304 900 -11104
rect 290 -11660 490 -11460
rect 1050 -12010 1250 -11810
<< metal2 >>
rect 1070 5680 1270 5689
rect 2835 5680 3025 5684
rect 1064 5480 1070 5680
rect 1270 5480 1276 5680
rect 2824 5675 3036 5680
rect 2824 5485 2835 5675
rect 3025 5485 3036 5675
rect 2824 5480 3036 5485
rect -740 1246 -540 1250
rect 1070 1246 1270 5480
rect 2830 1660 3030 5480
rect 2830 1460 6510 1660
rect -740 1046 1270 1246
rect 6310 1050 6510 1460
rect -546 -744 -540 -544
rect -340 -744 1090 -544
rect -146 -1104 -140 -904
rect 60 -1104 1090 -904
rect 290 -1274 490 -1268
rect 490 -1474 1090 -1274
rect 290 -1480 490 -1474
rect 698 -1624 898 -1618
rect 898 -1824 1090 -1624
rect 698 -1830 898 -1824
rect -740 -2614 -540 -2610
rect -740 -2814 1090 -2614
rect 6970 -2884 7170 -2880
rect -740 -3014 -540 -3010
rect -740 -3214 1090 -3014
rect 6510 -3084 7170 -2884
rect 6970 -3244 7170 -3240
rect 6504 -3444 7170 -3244
rect 6970 -3664 7170 -3660
rect 6504 -3864 7170 -3664
rect 6970 -4054 7170 -4050
rect 6510 -4254 7170 -4054
rect -740 -4274 -540 -4270
rect -740 -4474 1090 -4274
rect -740 -4684 -540 -4680
rect -740 -4884 1090 -4684
rect -740 -8380 -540 -8180
rect -340 -8184 -334 -8180
rect -340 -8380 1600 -8184
rect -740 -8384 1600 -8380
rect -130 -8804 70 -8798
rect 70 -9004 1600 -8804
rect -130 -9010 70 -9004
rect -740 -9314 -540 -9310
rect -740 -9514 1050 -9314
rect 1250 -9514 1600 -9314
rect -740 -9654 -540 -9650
rect -740 -9854 1600 -9654
rect -740 -10014 -540 -10010
rect 290 -10014 490 -10008
rect -740 -10214 290 -10014
rect 490 -10214 1600 -10014
rect 290 -10220 490 -10214
rect -740 -10404 -540 -10400
rect 6970 -10404 7170 -10396
rect -740 -10604 1600 -10404
rect 5650 -10604 7170 -10404
rect -740 -10744 -540 -10740
rect -740 -10944 290 -10744
rect 490 -10944 1600 -10744
rect 694 -11304 700 -11104
rect 900 -11304 1600 -11104
rect 284 -11660 290 -11460
rect 490 -11660 6650 -11460
rect 1050 -11810 1250 -11804
rect 1250 -12010 4880 -11810
rect 1050 -12016 1250 -12010
rect 4680 -14670 4880 -12010
rect 6450 -14670 6650 -11660
rect 4671 -14870 4680 -14670
rect 4880 -14870 4889 -14670
rect 6441 -14870 6450 -14670
rect 6650 -14870 6659 -14670
<< via2 >>
rect 1070 5480 1270 5680
rect 2835 5485 3025 5675
rect 4680 -14870 4880 -14670
rect 6450 -14870 6650 -14670
<< metal3 >>
rect 1065 5680 1275 5685
rect 1065 5475 1070 5680
rect 1270 5675 1275 5680
rect 2830 5679 3030 5680
rect 2825 5481 2831 5679
rect 3029 5481 3035 5679
rect 2830 5480 3030 5481
rect 1065 5469 1275 5475
rect 6445 -14665 6655 -14659
rect 4669 -14875 4675 -14665
rect 4875 -14670 4885 -14665
rect 4880 -14870 4885 -14670
rect 4875 -14875 4885 -14870
rect 6445 -14870 6450 -14865
rect 6650 -14870 6655 -14865
rect 6445 -14875 6655 -14870
<< via3 >>
rect 1070 5480 1270 5675
rect 1270 5480 1275 5675
rect 2831 5675 3029 5679
rect 2831 5485 2835 5675
rect 2835 5485 3025 5675
rect 3025 5485 3029 5675
rect 2831 5481 3029 5485
rect 1070 5475 1275 5480
rect 4675 -14670 4875 -14665
rect 4675 -14870 4680 -14670
rect 4680 -14870 4875 -14670
rect 4675 -14875 4875 -14870
rect 6445 -14670 6655 -14665
rect 6445 -14865 6450 -14670
rect 6450 -14865 6650 -14670
rect 6650 -14865 6655 -14670
<< metal4 >>
rect 1060 5675 1280 5680
rect 1060 5475 1070 5675
rect 1275 5475 1280 5675
rect 1060 5470 1280 5475
rect 2830 5679 3030 5680
rect 2830 5481 2831 5679
rect 3029 5481 3030 5679
rect 1070 -14530 1270 5470
rect 2830 -14540 3030 5481
rect 4675 -14664 4875 5410
rect 6450 -14664 6650 5410
rect 4674 -14665 4876 -14664
rect 4674 -14875 4675 -14665
rect 4875 -14875 4876 -14665
rect 6444 -14665 6656 -14664
rect 6444 -14865 6445 -14665
rect 6655 -14865 6656 -14665
rect 6444 -14866 6656 -14865
rect 4674 -14876 4876 -14875
use power_gating_ad  power_gating_ad_1
timestamp 1713788423
transform 1 0 760 0 1 -484
box -736 -8666 8950 3936
use power_gating_dd  power_gating_dd_0
timestamp 1713441137
transform 1 0 690 0 1 -5924
box 710 -5386 5190 -1514
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC3
timestamp 1713748097
transform 1 0 1296 0 1 -4550
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC4
timestamp 1713748097
transform 1 0 4916 0 1 -4550
box -1686 -9960 1686 9960
<< labels >>
flabel metal2 -740 1050 -540 1250 0 FreeSans 256 0 0 0 AVDD
port 6 nsew
flabel metal2 -740 -4470 -540 -4270 0 FreeSans 256 0 0 0 XIN
port 16 nsew
flabel metal2 -740 -4880 -540 -4680 0 FreeSans 256 0 0 0 AVSS
port 14 nsew
flabel metal2 -740 -9850 -540 -9650 0 FreeSans 256 0 0 0 SG_DVDD
port 5 nsew
flabel metal2 -740 -8380 -540 -8180 0 FreeSans 256 0 0 0 ENA
port 9 nsew
flabel metal2 -740 -10600 -540 -10400 0 FreeSans 256 0 0 0 SG_DVSS
port 10 nsew
flabel metal2 -740 -10210 -540 -10010 0 FreeSans 256 0 0 0 STDBY
port 12 nsew
flabel metal2 -740 -10940 -540 -10740 0 FreeSans 256 0 0 0 DVSS
port 15 nsew
flabel metal2 -740 -9510 -540 -9310 0 FreeSans 256 0 0 0 DVDD
port 3 nsew
flabel metal2 6970 -10596 7170 -10396 0 FreeSans 256 0 0 0 DOUT
port 1 nsew
flabel metal2 6970 -3860 7170 -3660 0 FreeSans 256 0 0 0 EG_AVSS
port 13 nsew
flabel metal2 6970 -3440 7170 -3240 0 FreeSans 256 0 0 0 EG_AVDD
port 8 nsew
flabel metal2 6970 -4250 7170 -4050 0 FreeSans 256 0 0 0 SG_AVSS
port 11 nsew
flabel metal2 6970 -3080 7170 -2880 0 FreeSans 256 0 0 0 SG_AVDD
port 2 nsew
flabel metal2 -740 -3210 -540 -3010 0 FreeSans 256 0 0 0 EG_IBIAS
port 4 nsew
flabel metal2 -740 -2810 -540 -2610 0 FreeSans 256 0 0 0 IBIAS
port 7 nsew
<< end >>
