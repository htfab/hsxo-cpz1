magic
tech sky130A
magscale 1 2
timestamp 1713748097
<< metal3 >>
rect -1686 9812 1686 9840
rect -1686 6788 1602 9812
rect 1666 6788 1686 9812
rect -1686 6760 1686 6788
rect -1686 6492 1686 6520
rect -1686 3468 1602 6492
rect 1666 3468 1686 6492
rect -1686 3440 1686 3468
rect -1686 3172 1686 3200
rect -1686 148 1602 3172
rect 1666 148 1686 3172
rect -1686 120 1686 148
rect -1686 -148 1686 -120
rect -1686 -3172 1602 -148
rect 1666 -3172 1686 -148
rect -1686 -3200 1686 -3172
rect -1686 -3468 1686 -3440
rect -1686 -6492 1602 -3468
rect 1666 -6492 1686 -3468
rect -1686 -6520 1686 -6492
rect -1686 -6788 1686 -6760
rect -1686 -9812 1602 -6788
rect 1666 -9812 1686 -6788
rect -1686 -9840 1686 -9812
<< via3 >>
rect 1602 6788 1666 9812
rect 1602 3468 1666 6492
rect 1602 148 1666 3172
rect 1602 -3172 1666 -148
rect 1602 -6492 1666 -3468
rect 1602 -9812 1666 -6788
<< mimcap >>
rect -1646 9760 1354 9800
rect -1646 6840 -1606 9760
rect 1314 6840 1354 9760
rect -1646 6800 1354 6840
rect -1646 6440 1354 6480
rect -1646 3520 -1606 6440
rect 1314 3520 1354 6440
rect -1646 3480 1354 3520
rect -1646 3120 1354 3160
rect -1646 200 -1606 3120
rect 1314 200 1354 3120
rect -1646 160 1354 200
rect -1646 -200 1354 -160
rect -1646 -3120 -1606 -200
rect 1314 -3120 1354 -200
rect -1646 -3160 1354 -3120
rect -1646 -3520 1354 -3480
rect -1646 -6440 -1606 -3520
rect 1314 -6440 1354 -3520
rect -1646 -6480 1354 -6440
rect -1646 -6840 1354 -6800
rect -1646 -9760 -1606 -6840
rect 1314 -9760 1354 -6840
rect -1646 -9800 1354 -9760
<< mimcapcontact >>
rect -1606 6840 1314 9760
rect -1606 3520 1314 6440
rect -1606 200 1314 3120
rect -1606 -3120 1314 -200
rect -1606 -6440 1314 -3520
rect -1606 -9760 1314 -6840
<< metal4 >>
rect -198 9761 -94 9960
rect 1582 9812 1686 9960
rect -1607 9760 1315 9761
rect -1607 6840 -1606 9760
rect 1314 6840 1315 9760
rect -1607 6839 1315 6840
rect -198 6441 -94 6839
rect 1582 6788 1602 9812
rect 1666 6788 1686 9812
rect 1582 6492 1686 6788
rect -1607 6440 1315 6441
rect -1607 3520 -1606 6440
rect 1314 3520 1315 6440
rect -1607 3519 1315 3520
rect -198 3121 -94 3519
rect 1582 3468 1602 6492
rect 1666 3468 1686 6492
rect 1582 3172 1686 3468
rect -1607 3120 1315 3121
rect -1607 200 -1606 3120
rect 1314 200 1315 3120
rect -1607 199 1315 200
rect -198 -199 -94 199
rect 1582 148 1602 3172
rect 1666 148 1686 3172
rect 1582 -148 1686 148
rect -1607 -200 1315 -199
rect -1607 -3120 -1606 -200
rect 1314 -3120 1315 -200
rect -1607 -3121 1315 -3120
rect -198 -3519 -94 -3121
rect 1582 -3172 1602 -148
rect 1666 -3172 1686 -148
rect 1582 -3468 1686 -3172
rect -1607 -3520 1315 -3519
rect -1607 -6440 -1606 -3520
rect 1314 -6440 1315 -3520
rect -1607 -6441 1315 -6440
rect -198 -6839 -94 -6441
rect 1582 -6492 1602 -3468
rect 1666 -6492 1686 -3468
rect 1582 -6788 1686 -6492
rect -1607 -6840 1315 -6839
rect -1607 -9760 -1606 -6840
rect 1314 -9760 1315 -6840
rect -1607 -9761 1315 -9760
rect -198 -9960 -94 -9761
rect 1582 -9812 1602 -6788
rect 1666 -9812 1686 -6788
rect 1582 -9960 1686 -9812
<< properties >>
string FIXED_BBOX -1686 6760 1394 9840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.0 l 15.0 val 461.4 carea 2.00 cperi 0.19 nx 1 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
