magic
tech sky130A
magscale 1 2
timestamp 1713441137
<< nwell >>
rect 1400 -3210 2070 -1720
rect 2490 -2360 3740 -1720
rect 1400 -4040 2100 -3210
<< pwell >>
rect 2500 -2980 3740 -2360
rect 3470 -4310 4160 -2980
rect 2820 -5130 3470 -4310
<< locali >>
rect 2092 -1744 2470 -1738
rect 3762 -1744 4140 -1738
rect 2086 -1812 2476 -1744
rect 2086 -1940 2160 -1812
rect 1310 -2140 2160 -1940
rect 2086 -2270 2160 -2140
rect 2402 -2270 2476 -1812
rect 3756 -1812 4146 -1744
rect 3756 -1940 3830 -1812
rect 3200 -1946 3830 -1940
rect 3200 -2134 3206 -1946
rect 3394 -2134 3830 -1946
rect 3200 -2140 3830 -2134
rect 2086 -2338 2476 -2270
rect 3756 -2270 3830 -2140
rect 4072 -2270 4146 -1812
rect 3756 -2338 4146 -2270
rect 2092 -2340 2470 -2338
rect 3762 -2340 4140 -2338
rect 2092 -2382 2470 -2380
rect 3762 -2382 4140 -2380
rect 2086 -2450 2476 -2382
rect 2086 -2890 2160 -2450
rect 2402 -2890 2476 -2450
rect 3756 -2450 4146 -2382
rect 3756 -2760 3830 -2450
rect 2086 -2958 2476 -2890
rect 3580 -2890 3830 -2760
rect 4072 -2890 4146 -2450
rect 3580 -2958 4146 -2890
rect 2092 -2964 2470 -2958
rect 3580 -2964 4140 -2958
rect 3580 -3026 3780 -2964
rect 3580 -3214 3586 -3026
rect 3774 -3214 3780 -3026
rect 3580 -3220 3780 -3214
rect 2122 -3234 2796 -3228
rect 2116 -3302 2802 -3234
rect 2116 -3390 2190 -3302
rect 1510 -3396 2190 -3390
rect 1694 -3584 2190 -3396
rect 1510 -3590 2190 -3584
rect 2116 -3960 2190 -3590
rect 2728 -3960 2802 -3302
rect 2116 -4028 2802 -3960
rect 2122 -4034 2796 -4028
rect 2124 -4332 2798 -4326
rect 3492 -4332 4166 -4326
rect 2118 -4400 2804 -4332
rect 2118 -5040 2192 -4400
rect 2730 -4760 2804 -4400
rect 3486 -4400 4172 -4332
rect 3486 -4760 3560 -4400
rect 2730 -4960 3560 -4760
rect 2730 -5040 2804 -4960
rect 2118 -5108 2804 -5040
rect 3486 -5040 3560 -4960
rect 4098 -4760 4172 -4400
rect 4098 -4766 4790 -4760
rect 4098 -4954 4596 -4766
rect 4784 -4954 4790 -4766
rect 4098 -4960 4790 -4954
rect 4098 -5040 4172 -4960
rect 3486 -5108 4172 -5040
rect 2124 -5114 2798 -5108
rect 3492 -5114 4166 -5108
<< viali >>
rect 1110 -2140 1310 -1940
rect 3206 -2134 3394 -1946
rect 3586 -3214 3774 -3026
rect 1506 -3584 1694 -3396
rect 4596 -4954 4784 -4766
<< metal1 >>
rect 1494 -1720 1500 -1520
rect 1700 -1720 1706 -1520
rect 1104 -1940 1316 -1928
rect 1104 -2140 1110 -1940
rect 1310 -2140 1316 -1940
rect 1104 -2152 1316 -2140
rect 1110 -3390 1310 -2152
rect 1500 -2880 1700 -1720
rect 3200 -1940 3400 -1934
rect 3194 -2140 3200 -1940
rect 3400 -2140 3406 -1940
rect 2804 -2460 2810 -2260
rect 3010 -2460 3016 -2260
rect 1494 -3080 1500 -2880
rect 1700 -3080 1706 -2880
rect 2810 -3190 3010 -2460
rect 1500 -3390 1700 -3384
rect 1104 -3590 1110 -3390
rect 1310 -3590 1316 -3390
rect 1500 -3596 1700 -3590
rect 1900 -3390 3010 -3190
rect 1900 -3870 2100 -3390
rect 2240 -3443 2294 -3433
rect 2240 -3597 2294 -3587
rect 2432 -3443 2486 -3433
rect 2432 -3597 2486 -3587
rect 2624 -3443 2678 -3433
rect 2624 -3597 2678 -3587
rect 2336 -3675 2390 -3665
rect 2336 -3829 2390 -3819
rect 2528 -3675 2582 -3665
rect 2528 -3829 2582 -3819
rect 2810 -3870 3010 -3390
rect 3200 -3390 3400 -2140
rect 4320 -2260 4520 -2254
rect 3574 -3220 3580 -3020
rect 3780 -3220 3786 -3020
rect 4320 -3040 4520 -2460
rect 3200 -3596 3400 -3590
rect 4120 -3240 4520 -3040
rect 1500 -4070 3470 -3870
rect 1500 -4090 1700 -4070
rect 2812 -4290 3012 -4284
rect 1500 -4296 1700 -4290
rect 1902 -4490 2812 -4290
rect 1902 -4960 2102 -4490
rect 2242 -4532 2296 -4522
rect 2242 -4686 2296 -4676
rect 2434 -4532 2488 -4522
rect 2434 -4686 2488 -4676
rect 2626 -4532 2680 -4522
rect 2626 -4686 2680 -4676
rect 2338 -4764 2392 -4754
rect 2338 -4918 2392 -4908
rect 2530 -4764 2584 -4754
rect 2530 -4918 2584 -4908
rect 2812 -4960 3012 -4490
rect 1500 -5160 3012 -4960
rect 3270 -4290 3470 -4070
rect 4120 -3970 4320 -3240
rect 4584 -3660 4590 -3460
rect 4790 -3660 4796 -3460
rect 4120 -4176 4320 -4170
rect 3270 -4490 4390 -4290
rect 3270 -4950 3470 -4490
rect 3610 -4532 3664 -4522
rect 3610 -4686 3664 -4676
rect 3802 -4532 3856 -4522
rect 3802 -4686 3856 -4676
rect 3994 -4532 4048 -4522
rect 3994 -4686 4048 -4676
rect 3706 -4764 3760 -4754
rect 3706 -4918 3760 -4908
rect 3898 -4764 3952 -4754
rect 3898 -4918 3952 -4908
rect 4190 -4950 4390 -4490
rect 3270 -5160 4390 -4950
rect 4590 -4760 4790 -3660
rect 4590 -4966 4790 -4960
rect 1500 -5180 1700 -5160
rect 1500 -5386 1700 -5380
<< via1 >>
rect 1500 -1720 1700 -1520
rect 3200 -1946 3400 -1940
rect 3200 -2134 3206 -1946
rect 3206 -2134 3394 -1946
rect 3394 -2134 3400 -1946
rect 3200 -2140 3400 -2134
rect 2810 -2460 3010 -2260
rect 1500 -3080 1700 -2880
rect 1110 -3590 1310 -3390
rect 1500 -3396 1700 -3390
rect 1500 -3584 1506 -3396
rect 1506 -3584 1694 -3396
rect 1694 -3584 1700 -3396
rect 1500 -3590 1700 -3584
rect 2240 -3587 2294 -3443
rect 2432 -3587 2486 -3443
rect 2624 -3587 2678 -3443
rect 2336 -3819 2390 -3675
rect 2528 -3819 2582 -3675
rect 4320 -2460 4520 -2260
rect 3580 -3026 3780 -3020
rect 3580 -3214 3586 -3026
rect 3586 -3214 3774 -3026
rect 3774 -3214 3780 -3026
rect 3580 -3220 3780 -3214
rect 3200 -3590 3400 -3390
rect 1500 -4290 1700 -4090
rect 2812 -4490 3012 -4290
rect 2242 -4676 2296 -4532
rect 2434 -4676 2488 -4532
rect 2626 -4676 2680 -4532
rect 2338 -4908 2392 -4764
rect 2530 -4908 2584 -4764
rect 4590 -3660 4790 -3460
rect 4120 -4170 4320 -3970
rect 3610 -4676 3664 -4532
rect 3802 -4676 3856 -4532
rect 3994 -4676 4048 -4532
rect 3706 -4908 3760 -4764
rect 3898 -4908 3952 -4764
rect 4590 -4766 4790 -4760
rect 4590 -4954 4596 -4766
rect 4596 -4954 4784 -4766
rect 4784 -4954 4790 -4766
rect 4590 -4960 4790 -4954
rect 1500 -5380 1700 -5180
<< metal2 >>
rect 1500 -1520 1700 -1514
rect 1700 -1720 2650 -1520
rect 1500 -1726 1700 -1720
rect 1910 -2140 2110 -1940
rect 710 -2460 2110 -2260
rect 2450 -2460 2650 -1720
rect 3200 -1940 3400 -1934
rect 3400 -2140 3770 -1940
rect 3200 -2146 3400 -2140
rect 2810 -2260 3010 -2254
rect 3010 -2460 3780 -2260
rect 4120 -2460 4320 -2260
rect 4520 -2460 4526 -2260
rect 2810 -2466 3010 -2460
rect 1500 -2880 1700 -2874
rect 710 -3080 1500 -2880
rect 1500 -3086 1700 -3080
rect 1910 -3020 2110 -2570
rect 2810 -2770 3780 -2570
rect 2810 -3020 3010 -2770
rect 1910 -3220 3010 -3020
rect 3580 -3020 3780 -2770
rect 1110 -3390 1310 -3384
rect 710 -3590 1110 -3390
rect 1310 -3590 1500 -3390
rect 1700 -3443 3200 -3390
rect 1700 -3587 2240 -3443
rect 2294 -3587 2432 -3443
rect 2486 -3587 2624 -3443
rect 2678 -3587 3200 -3443
rect 1700 -3590 3200 -3587
rect 3400 -3590 3406 -3390
rect 3580 -3460 3780 -3220
rect 4590 -3460 4790 -3454
rect 1110 -3596 1310 -3590
rect 3580 -3660 4590 -3460
rect 4590 -3666 4790 -3660
rect 1500 -3675 2680 -3670
rect 1500 -3730 2336 -3675
rect 710 -3819 2336 -3730
rect 2390 -3819 2528 -3675
rect 2582 -3819 2680 -3675
rect 710 -3870 2680 -3819
rect 710 -3930 1700 -3870
rect 710 -4290 1500 -4090
rect 1700 -4290 1706 -4090
rect 2812 -4170 4120 -3970
rect 4320 -4170 4326 -3970
rect 2812 -4290 3012 -4170
rect 710 -4532 2690 -4480
rect 2806 -4490 2812 -4290
rect 3012 -4490 3018 -4290
rect 710 -4676 2242 -4532
rect 2296 -4676 2434 -4532
rect 2488 -4676 2626 -4532
rect 2680 -4676 2690 -4532
rect 710 -4680 2690 -4676
rect 3600 -4532 5190 -4480
rect 3600 -4676 3610 -4532
rect 3664 -4676 3802 -4532
rect 3856 -4676 3994 -4532
rect 4048 -4676 5190 -4532
rect 3600 -4680 5190 -4676
rect 1500 -4764 4590 -4760
rect 1500 -4820 2338 -4764
rect 710 -4908 2338 -4820
rect 2392 -4908 2530 -4764
rect 2584 -4908 3706 -4764
rect 3760 -4908 3898 -4764
rect 3952 -4908 4590 -4764
rect 710 -4960 4590 -4908
rect 4790 -4960 4796 -4760
rect 710 -5020 1700 -4960
rect 710 -5380 1500 -5180
rect 1700 -5380 1706 -5180
use level_shifter_dd  level_shifter_dd_0
timestamp 1713441137
transform 1 0 1690 0 1 -1070
box 220 -1910 960 -652
use level_shifter_dd  level_shifter_dd_1
timestamp 1713441137
transform 1 0 3360 0 1 -1070
box 220 -1910 960 -652
use sky130_fd_pr__nfet_01v8_F5PS5H  XM4
timestamp 1713252812
transform 1 0 3829 0 1 -4720
box -359 -410 359 410
use sky130_fd_pr__nfet_01v8_F5PS5H  XM18
timestamp 1713252812
transform 1 0 2461 0 1 -4720
box -359 -410 359 410
use sky130_fd_pr__pfet_01v8_XG6UDL  XM27
timestamp 1713252812
transform 1 0 2459 0 1 -3631
box -359 -419 359 419
<< labels >>
flabel metal2 4990 -4680 5190 -4480 0 FreeSans 256 0 0 0 DOUT
port 8 nsew
flabel metal2 710 -2460 910 -2260 0 FreeSans 256 0 0 0 ENA
port 2 nsew
flabel metal2 710 -3080 910 -2880 0 FreeSans 256 0 0 0 ENA_B
port 3 nsew
flabel metal2 710 -3590 910 -3390 0 FreeSans 256 0 0 0 DVDD
port 1 nsew
flabel metal2 710 -4290 910 -4090 0 FreeSans 256 0 0 0 STDBY
port 4 nsew
flabel metal2 710 -4680 910 -4480 0 FreeSans 256 0 0 0 SG_DVSS
port 6 nsew
flabel metal2 710 -5380 910 -5180 0 FreeSans 256 0 0 0 STDBY_B
port 5 nsew
flabel metal2 710 -3930 910 -3730 0 FreeSans 256 0 0 0 SG_DVDD
port 7 nsew
flabel metal2 710 -5020 910 -4820 0 FreeSans 256 0 0 0 DVSS
port 0 nsew
<< end >>
