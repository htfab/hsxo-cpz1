magic
tech sky130A
magscale 1 2
timestamp 1713249940
<< error_s >>
rect 440 -4920 960 -4320
rect 1040 -5020 6710 -3760
rect 6760 -5020 7310 -4320
<< dnwell >>
rect 960 -4920 6760 1550
rect 960 -5020 1040 -4920
rect 6710 -5020 6760 -4920
rect 960 -5240 6760 -5020
rect 2110 -11280 5650 -7180
<< nwell >>
rect 850 930 6870 1660
rect 850 740 1570 930
rect 850 -2614 1370 740
rect 5530 130 6870 930
rect 850 -2814 1720 -2614
rect 850 -3160 1370 -2814
rect 850 -3360 4500 -3160
rect 850 -4920 1166 -3360
rect 6554 -4920 6870 130
rect 850 -5350 6870 -4920
rect 2030 -7386 5730 -7100
rect 2030 -11074 2316 -7386
rect 5444 -11074 5730 -7386
rect 2030 -11360 5730 -11074
<< nsubdiff >>
rect 2067 -7157 5693 -7137
rect 2067 -7191 2147 -7157
rect 5613 -7191 5693 -7157
rect 2067 -7211 5693 -7191
rect 2067 -7217 2141 -7211
rect 2067 -11243 2087 -7217
rect 2121 -11243 2141 -7217
rect 2067 -11249 2141 -11243
rect 5619 -7217 5693 -7211
rect 5619 -11243 5639 -7217
rect 5673 -11243 5693 -7217
rect 5619 -11249 5693 -11243
rect 2067 -11269 5693 -11249
rect 2067 -11303 2147 -11269
rect 5613 -11303 5693 -11269
rect 2067 -11323 5693 -11303
<< mvnsubdiff >>
rect 917 1573 6803 1593
rect 917 1539 997 1573
rect 6723 1539 6803 1573
rect 917 1519 6803 1539
rect 917 1513 991 1519
rect 917 -5203 937 1513
rect 971 -5203 991 1513
rect 917 -5209 991 -5203
rect 6729 1513 6803 1519
rect 6729 -5203 6749 1513
rect 6783 -5203 6803 1513
rect 6729 -5209 6803 -5203
rect 917 -5229 6803 -5209
rect 917 -5263 997 -5229
rect 6723 -5263 6803 -5229
rect 917 -5283 6803 -5263
<< nsubdiffcont >>
rect 2147 -7191 5613 -7157
rect 2087 -11243 2121 -7217
rect 5639 -11243 5673 -7217
rect 2147 -11303 5613 -11269
<< mvnsubdiffcont >>
rect 997 1539 6723 1573
rect 937 -5203 971 1513
rect 6749 -5203 6783 1513
rect 997 -5263 6723 -5229
<< locali >>
rect 937 1539 997 1573
rect 6723 1539 6783 1573
rect 937 1513 971 1539
rect 937 -5229 971 -5203
rect 6749 1513 6783 1539
rect 6749 -5229 6783 -5203
rect 937 -5263 997 -5229
rect 6723 -5263 6783 -5229
rect 2087 -7191 2147 -7157
rect 5613 -7191 5673 -7157
rect 2087 -7217 2121 -7191
rect 2087 -11269 2121 -11243
rect 5639 -7217 5673 -7191
rect 5639 -11269 5673 -11243
rect 2087 -11303 2147 -11269
rect 5613 -11303 5673 -11269
<< metal2 >>
rect 520 1046 1740 1246
rect -1770 10 -1570 210
rect -1770 -390 -1570 -190
rect -1770 -790 -1570 -590
rect -1770 -1190 -1570 -990
rect -1770 -1590 -1570 -1390
rect -1770 -1990 -1570 -1790
rect -1770 -2390 -1570 -2190
rect -1770 -2790 -1570 -2590
rect 3900 -2850 4100 -1719
rect -1770 -3190 -1570 -2990
rect -1770 -3590 -1570 -3390
rect -1770 -3990 -1570 -3790
rect -1770 -4390 -1570 -4190
rect -1770 -4790 -1570 -4590
rect -1770 -5190 -1570 -4990
rect -1770 -5590 -1570 -5390
use power_gating_ad  power_gating_ad_0
timestamp 1713249912
transform 1 0 960 0 1 -484
box 130 -4406 5950 1736
use power_gating_dd  power_gating_dd_0
timestamp 1713242883
transform 1 0 690 0 1 -5924
box 1110 -5386 5190 -1720
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC3
timestamp 1713241921
transform 1 0 9176 0 1 -12920
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC4
timestamp 1713241921
transform 1 0 13586 0 1 -12800
box -1686 -9960 1686 9960
<< labels >>
flabel metal2 -1770 10 -1570 210 0 FreeSans 256 0 0 0 DOUT
port 0 nsew
flabel metal2 -1770 -390 -1570 -190 0 FreeSans 256 0 0 0 SG_AVDD
port 1 nsew
flabel metal2 -1770 -790 -1570 -590 0 FreeSans 256 0 0 0 DVDD
port 2 nsew
flabel metal2 -1770 -1190 -1570 -990 0 FreeSans 256 0 0 0 EG_IBIAS
port 3 nsew
flabel metal2 -1770 -1590 -1570 -1390 0 FreeSans 256 0 0 0 SG_DVDD
port 4 nsew
flabel metal2 -1770 -1990 -1570 -1790 0 FreeSans 256 0 0 0 AVDD
port 5 nsew
flabel metal2 -1770 -2390 -1570 -2190 0 FreeSans 256 0 0 0 IBIAS
port 6 nsew
flabel metal2 -1770 -2790 -1570 -2590 0 FreeSans 256 0 0 0 EG_AVDD
port 7 nsew
flabel metal2 -1770 -3190 -1570 -2990 0 FreeSans 256 0 0 0 ENA
port 8 nsew
flabel metal2 -1770 -3590 -1570 -3390 0 FreeSans 256 0 0 0 SG_DVSS
port 9 nsew
flabel metal2 -1770 -3990 -1570 -3790 0 FreeSans 256 0 0 0 SG_AVSS
port 10 nsew
flabel metal2 -1770 -4390 -1570 -4190 0 FreeSans 256 0 0 0 STDBY
port 11 nsew
flabel metal2 -1770 -4790 -1570 -4590 0 FreeSans 256 0 0 0 EG_AVSS
port 12 nsew
flabel metal2 -1770 -5190 -1570 -4990 0 FreeSans 256 0 0 0 AVSS
port 13 nsew
flabel metal2 -1770 -5590 -1570 -5390 0 FreeSans 256 0 0 0 DVSS
port 14 nsew
<< end >>
