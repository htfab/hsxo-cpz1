magic
tech sky130A
magscale 1 2
timestamp 1713242186
<< dnwell >>
rect 60 -3010 1840 780
rect 3550 -3050 6100 1030
<< nwell >>
rect -20 -1490 1920 860
rect -20 -2804 266 -1490
rect 1634 -2804 1920 -1490
rect -20 -3090 1920 -2804
rect 3440 -1390 6210 1140
rect 3440 -2844 3756 -1390
rect 5894 -2844 6210 -1390
rect 3440 -3160 6210 -2844
<< psubdiff >>
rect 740 -2170 1140 -2146
rect 740 -2594 1140 -2570
<< nsubdiff >>
rect 17 803 1883 823
rect 17 769 97 803
rect 1803 769 1883 803
rect 17 749 1883 769
rect 17 743 91 749
rect 17 -2973 37 743
rect 71 -2973 91 743
rect 1809 743 1883 749
rect 750 80 1150 104
rect 750 -344 1150 -320
rect 17 -2979 91 -2973
rect 1809 -2973 1829 743
rect 1863 -2973 1883 743
rect 1809 -2979 1883 -2973
rect 17 -2999 1883 -2979
rect 17 -3033 97 -2999
rect 1803 -3033 1883 -2999
rect 17 -3053 1883 -3033
<< mvpsubdiff >>
rect 4580 -2220 4980 -2196
rect 4580 -2644 4980 -2620
<< mvnsubdiff >>
rect 3507 1053 6143 1073
rect 3507 1019 3587 1053
rect 6063 1019 6143 1053
rect 3507 999 6143 1019
rect 3507 993 3581 999
rect 3507 -3013 3527 993
rect 3561 -3013 3581 993
rect 6069 993 6143 999
rect 4280 300 4680 324
rect 4280 -124 4680 -100
rect 3507 -3019 3581 -3013
rect 6069 -3013 6089 993
rect 6123 -3013 6143 993
rect 6069 -3019 6143 -3013
rect 3507 -3039 6143 -3019
rect 3507 -3073 3587 -3039
rect 6063 -3073 6143 -3039
rect 3507 -3093 6143 -3073
<< psubdiffcont >>
rect 740 -2570 1140 -2170
<< nsubdiffcont >>
rect 97 769 1803 803
rect 37 -2973 71 743
rect 750 -320 1150 80
rect 1829 -2973 1863 743
rect 97 -3033 1803 -2999
<< mvpsubdiffcont >>
rect 4580 -2620 4980 -2220
<< mvnsubdiffcont >>
rect 3587 1019 6063 1053
rect 3527 -3013 3561 993
rect 4280 -100 4680 300
rect 6089 -3013 6123 993
rect 3587 -3073 6063 -3039
<< locali >>
rect 3527 1019 3587 1053
rect 6063 1019 6123 1053
rect 3527 993 3561 1019
rect 37 769 97 803
rect 1803 769 1863 803
rect 37 743 71 769
rect 1829 743 1863 769
rect 750 80 1150 96
rect 750 -336 1150 -320
rect 740 -2170 1140 -2154
rect 740 -2586 1140 -2570
rect 37 -2999 71 -2973
rect 1829 -2999 1863 -2973
rect 37 -3033 97 -2999
rect 1803 -3033 1863 -2999
rect 6089 993 6123 1019
rect 4280 300 4680 316
rect 4280 -116 4680 -100
rect 4580 -2220 4980 -2204
rect 4580 -2636 4980 -2620
rect 3527 -3039 3561 -3013
rect 6089 -3039 6123 -3013
rect 3527 -3073 3587 -3039
rect 6063 -3073 6123 -3039
<< viali >>
rect 4686 -2514 4874 -2326
<< metal1 >>
rect 4380 200 4580 206
rect 850 -10 1050 -4
rect 4380 -6 4580 0
rect 850 -216 1050 -210
rect 2490 -1390 2690 -1384
rect 194 -1590 200 -1390
rect 400 -1590 406 -1390
rect 200 -2770 400 -1590
rect 1870 -2070 2070 -2064
rect 840 -2270 1040 -2264
rect 840 -2476 1040 -2470
rect 200 -2976 400 -2970
rect 1870 -2770 2070 -2270
rect 2490 -2770 2690 -1590
rect 4674 -2520 4680 -2320
rect 4880 -2520 4886 -2320
rect 2484 -2970 2490 -2770
rect 2690 -2970 2696 -2770
rect 1870 -2976 2070 -2970
<< via1 >>
rect 4380 0 4580 200
rect 850 -210 1050 -10
rect 200 -1590 400 -1390
rect 2490 -1590 2690 -1390
rect 840 -2470 1040 -2270
rect 1870 -2270 2070 -2070
rect 200 -2970 400 -2770
rect 4680 -2326 4880 -2320
rect 4680 -2514 4686 -2326
rect 4686 -2514 4874 -2326
rect 4874 -2514 4880 -2326
rect 4680 -2520 4880 -2514
rect 1870 -2970 2070 -2770
rect 2490 -2970 2690 -2770
<< metal2 >>
rect 4374 0 4380 200
rect 4580 0 4880 200
rect 590 -210 850 -10
rect 1050 -210 1056 -10
rect 590 -1270 790 -210
rect 4680 -710 4880 0
rect 200 -1390 400 -1384
rect 400 -1590 790 -1390
rect 1130 -1590 2490 -1390
rect 2690 -1590 2696 -1390
rect 4070 -1480 4270 -1280
rect 5300 -1480 5500 -1280
rect 200 -1596 400 -1590
rect 590 -2270 790 -1700
rect 1864 -2270 1870 -2070
rect 2070 -2270 4580 -2070
rect 590 -2470 840 -2270
rect 1040 -2470 1046 -2270
rect 4680 -2320 4880 -2070
rect 4680 -2526 4880 -2520
rect 2490 -2770 2690 -2764
rect 4990 -2770 5190 -2070
rect 194 -2970 200 -2770
rect 400 -2970 1870 -2770
rect 2070 -2970 2076 -2770
rect 2690 -2970 5190 -2770
rect 2490 -2976 2690 -2970
use level_shifter_ad  level_shifter_ad_0
timestamp 1713241808
transform 1 0 3190 0 1 -300
box 880 -1970 2310 -210
use level_shifter_dd  level_shifter_dd_1
timestamp 1713242186
transform 1 0 370 0 1 -200
box 220 -1910 960 -652
<< labels >>
flabel metal2 590 -1270 790 -1070 0 FreeSans 256 0 0 0 DVDD
port 2 nsew
flabel metal2 590 -1900 790 -1700 0 FreeSans 256 0 0 0 DVSS
port 6 nsew
flabel metal2 590 -1590 790 -1390 0 FreeSans 256 0 0 0 LO
port 3 nsew
flabel metal2 1130 -1590 1330 -1390 0 FreeSans 256 0 0 0 LO_B
port 1 nsew
flabel metal2 4680 -710 4880 -510 0 FreeSans 256 0 0 0 AVDD
port 0 nsew
flabel metal2 4070 -1480 4270 -1280 0 FreeSans 256 0 0 0 HI_B
port 7 nsew
flabel metal2 4990 -2270 5190 -2070 0 FreeSans 256 0 0 0 LO_B
port 1 nsew
flabel metal2 4680 -2270 4880 -2070 0 FreeSans 256 0 0 0 AVSS
port 5 nsew
flabel metal2 5300 -1480 5500 -1280 0 FreeSans 256 0 0 0 HI
port 4 nsew
flabel metal2 4380 -2270 4580 -2070 0 FreeSans 256 0 0 0 LO
port 3 nsew
<< end >>
