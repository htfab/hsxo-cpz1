magic
tech sky130A
magscale 1 2
timestamp 1713782160
<< nwell >>
rect -200 2610 5370 2620
rect -200 1820 1120 2610
rect 2340 1820 4140 2610
rect 5360 1820 5370 2610
rect -200 -1860 980 1820
rect -200 -2870 5630 -1860
<< pwell >>
rect 1700 1050 1760 1770
rect 2320 1050 4160 1770
rect 4730 1050 4780 1770
rect 5330 1050 6110 1770
rect 1290 -6960 2410 -6830
rect 1290 -7330 1630 -6960
rect 1970 -7304 1990 -7300
rect 1970 -7324 1992 -7304
rect 2000 -7330 2410 -6960
rect 1290 -7460 2410 -7330
rect 3440 -7510 4610 -6610
rect 5640 -7520 6110 1050
<< locali >>
rect 1630 2924 1830 2930
rect 1630 2736 1636 2924
rect 1824 2736 1830 2924
rect 1630 2556 1830 2736
rect 4650 2924 4850 2930
rect 4650 2736 4656 2924
rect 4844 2736 4850 2924
rect 4650 2556 4850 2736
rect 1184 2550 2282 2556
rect 4204 2550 5302 2556
rect 1178 2482 2288 2550
rect 1178 1952 1252 2482
rect 1604 2350 1862 2482
rect 1604 1952 1678 2350
rect 1178 1884 1678 1952
rect 1788 1952 1862 2350
rect 2214 1952 2288 2482
rect 1788 1884 2288 1952
rect 4198 2482 5308 2550
rect 4198 1952 4272 2482
rect 4624 2350 4882 2482
rect 4624 1952 4698 2350
rect 4198 1884 4698 1952
rect 4808 1952 4882 2350
rect 5234 1952 5308 2482
rect 4808 1884 5308 1952
rect 1184 1878 1672 1884
rect 1794 1878 2282 1884
rect 4204 1878 4692 1884
rect 4814 1878 5302 1884
rect 1184 1734 1672 1738
rect 1794 1734 2282 1738
rect 1184 1732 2282 1734
rect 4204 1732 4692 1738
rect 4814 1732 5302 1738
rect 1178 1664 2288 1732
rect 1178 1152 1252 1664
rect 1604 1546 1862 1664
rect 1604 1152 1678 1546
rect 1178 1084 1678 1152
rect 1788 1152 1862 1546
rect 2214 1152 2288 1664
rect 1788 1084 2288 1152
rect 4198 1664 4698 1732
rect 4198 1152 4272 1664
rect 4624 1280 4698 1664
rect 4808 1664 5308 1732
rect 4808 1280 4882 1664
rect 4624 1152 4882 1280
rect 5234 1152 5308 1664
rect 4198 1084 5308 1152
rect 1184 1078 1672 1084
rect 1794 1078 2282 1084
rect 4204 1078 5302 1084
rect 4650 774 4850 1078
rect 4650 586 4656 774
rect 4844 586 4850 774
rect 4650 580 4850 586
rect 2860 -1724 2866 -1530
rect 3654 -1724 3660 -1680
rect 2860 -1920 3660 -1724
rect 1958 -1924 2482 -1920
rect 2760 -1924 4640 -1920
rect 1054 -1930 5566 -1924
rect 1048 -1998 5572 -1930
rect 1048 -2728 1122 -1998
rect 1948 -2125 2502 -1998
rect 1948 -2728 2022 -2125
rect 1048 -2730 2022 -2728
rect 570 -2796 2022 -2730
rect 2428 -2728 2502 -2125
rect 3328 -2120 4672 -1998
rect 3328 -2728 3402 -2120
rect 2428 -2796 3402 -2728
rect 4598 -2728 4672 -2120
rect 5498 -2728 5572 -1998
rect 4598 -2796 5572 -2728
rect 570 -2802 2016 -2796
rect 2434 -2802 3396 -2796
rect 4604 -2802 5566 -2796
rect 570 -2880 1370 -2802
rect 570 -3060 590 -2880
rect 1350 -3060 1370 -2880
rect 570 -3070 1370 -3060
rect 2444 -6638 3406 -6632
rect 4644 -6638 5606 -6632
rect 2438 -6706 3412 -6638
rect 565 -6750 1381 -6739
rect 565 -6830 580 -6750
rect 660 -6830 1290 -6750
rect 1370 -6830 1381 -6750
rect 565 -6840 1381 -6830
rect 565 -7450 670 -6840
rect 775 -6950 1171 -6949
rect 775 -7040 890 -6950
rect 1050 -7040 1171 -6950
rect 775 -7049 1171 -7040
rect 775 -7245 875 -7049
rect 1071 -7245 1171 -7049
rect 775 -7345 1171 -7245
rect 1280 -7450 1381 -6840
rect 1610 -6960 2014 -6945
rect 1610 -7030 1620 -6960
rect 1690 -7030 1930 -6960
rect 2000 -7030 2014 -6960
rect 1610 -7045 2014 -7030
rect 1610 -7249 1712 -7045
rect 1914 -7249 2014 -7045
rect 1610 -7270 2014 -7249
rect 1610 -7340 1620 -7270
rect 1690 -7340 1930 -7270
rect 2000 -7340 2014 -7270
rect 1610 -7349 2014 -7340
rect 565 -7460 1381 -7450
rect 2438 -7418 2512 -6706
rect 3338 -7295 3412 -6706
rect 4638 -6706 5612 -6638
rect 4638 -7295 4712 -6706
rect 3338 -7418 4712 -7295
rect 5538 -7418 5612 -6706
rect 2438 -7460 5612 -7418
rect 565 -7540 580 -7460
rect 660 -7540 1290 -7460
rect 1370 -7540 1381 -7460
rect 565 -7555 1381 -7540
rect 1920 -7466 5612 -7460
rect 1920 -7654 1926 -7466
rect 2114 -7486 5612 -7466
rect 2114 -7492 5606 -7486
rect 2114 -7654 2490 -7492
rect 3360 -7500 4692 -7492
rect 1920 -7660 2490 -7654
<< viali >>
rect 1636 2736 1824 2924
rect 4656 2736 4844 2924
rect 4656 586 4844 774
rect 2866 -1724 3654 -936
rect 590 -3060 1350 -2880
rect 580 -6830 660 -6750
rect 1290 -6830 1370 -6750
rect 890 -7040 1050 -6950
rect 1620 -7030 1690 -6960
rect 1930 -7030 2000 -6960
rect 1620 -7340 1690 -7270
rect 1930 -7340 2000 -7270
rect 580 -7540 660 -7460
rect 1290 -7540 1370 -7460
rect 1926 -7654 2114 -7466
<< metal1 >>
rect -270 3530 530 3536
rect 6350 3530 7150 3536
rect -276 2730 -270 2930
rect 1630 2930 1830 2936
rect 1624 2730 1630 2930
rect 1830 2730 1836 2930
rect 2854 2730 2860 3530
rect 3660 2730 3666 3530
rect 4650 2930 4850 2936
rect 4644 2730 4650 2930
rect 4850 2730 4856 2930
rect -270 -2870 530 2730
rect 1630 2724 1830 2730
rect 722 1727 728 1932
rect 933 1727 939 1932
rect 2300 1730 2330 1930
rect 2530 1730 2600 1930
rect 728 -1920 933 1727
rect 1934 940 1940 1140
rect 2140 940 2146 1140
rect 1940 780 2140 940
rect 1104 580 1110 780
rect 1310 580 2140 780
rect 2400 -928 2600 1730
rect 2112 -1133 2118 -928
rect 2323 -1133 2600 -928
rect 2860 -930 3660 2730
rect 4650 2724 4850 2730
rect 3918 1930 4103 1932
rect 5510 1930 5710 1936
rect 3918 1730 3960 1930
rect 4160 1730 4190 1930
rect 5505 1730 5510 1902
rect 3918 -928 4123 1730
rect 4344 940 4350 1140
rect 4550 940 4556 1140
rect 4954 940 4960 1140
rect 5160 940 5166 1140
rect 4350 -190 4550 940
rect 4650 780 4850 786
rect 4650 574 4850 580
rect 4344 -390 4350 -190
rect 4550 -390 4556 -190
rect 4960 -540 5160 940
rect 4960 -746 5160 -740
rect 3912 -1133 3918 -928
rect 4123 -1133 4129 -928
rect 2860 -1736 3660 -1730
rect 5505 -1920 5710 1730
rect 6350 780 7150 2730
rect 6344 -20 6350 780
rect 7150 -20 7156 780
rect 728 -2122 3540 -1920
rect 910 -2125 3540 -2122
rect 910 -2605 1115 -2125
rect 1192 -2175 1246 -2165
rect 1192 -2329 1246 -2319
rect 1508 -2175 1562 -2165
rect 1508 -2329 1562 -2319
rect 1824 -2175 1878 -2165
rect 1824 -2329 1878 -2319
rect 1350 -2407 1404 -2397
rect 1350 -2561 1404 -2551
rect 1666 -2407 1720 -2397
rect 1666 -2561 1720 -2551
rect 1955 -2605 2160 -2125
rect 910 -2810 2160 -2605
rect 2290 -2605 2495 -2125
rect 2572 -2175 2626 -2165
rect 2572 -2329 2626 -2319
rect 2888 -2175 2942 -2165
rect 2888 -2329 2942 -2319
rect 3204 -2175 3258 -2165
rect 3204 -2329 3258 -2319
rect 2730 -2407 2784 -2397
rect 2730 -2561 2784 -2551
rect 3046 -2407 3100 -2397
rect 3046 -2561 3100 -2551
rect 3335 -2605 3540 -2125
rect 2290 -2810 3540 -2605
rect 4460 -2125 5710 -1920
rect 4460 -2605 4665 -2125
rect 4742 -2175 4796 -2165
rect 4742 -2329 4796 -2319
rect 5058 -2175 5112 -2165
rect 5058 -2329 5112 -2319
rect 5374 -2175 5428 -2165
rect 5374 -2329 5428 -2319
rect 4900 -2407 4954 -2397
rect 4900 -2561 4954 -2551
rect 5216 -2407 5270 -2397
rect 5216 -2561 5270 -2551
rect 5505 -2605 5710 -2125
rect 4460 -2810 5710 -2605
rect 5937 -928 6142 -922
rect -270 -2880 1370 -2870
rect -270 -3060 590 -2880
rect 1350 -3060 1370 -2880
rect -270 -3870 1370 -3060
rect 570 -6460 1370 -3870
rect 515 -6750 715 -6700
rect 515 -6830 580 -6750
rect 660 -6830 715 -6750
rect 515 -7405 715 -6830
rect 871 -6950 1071 -6460
rect 871 -7040 890 -6950
rect 1050 -7040 1071 -6950
rect 871 -7050 1071 -7040
rect 1231 -6750 1431 -6690
rect 2112 -6703 2118 -6498
rect 2323 -6620 2495 -6498
rect 5937 -6620 6142 -1133
rect 2323 -6703 3540 -6620
rect 1231 -6830 1290 -6750
rect 1370 -6830 1431 -6750
rect 900 -7090 1040 -7080
rect 900 -7210 910 -7090
rect 1030 -7210 1040 -7090
rect 900 -7220 1040 -7210
rect 1231 -7260 1431 -6830
rect 2290 -6825 3540 -6703
rect 1500 -6960 2120 -6840
rect 1500 -7030 1620 -6960
rect 1690 -7030 1930 -6960
rect 2000 -7030 2120 -6960
rect 1500 -7040 2120 -7030
rect 1500 -7260 1700 -7040
rect 1740 -7090 1880 -7080
rect 1740 -7210 1750 -7090
rect 1870 -7210 1880 -7090
rect 1740 -7220 1880 -7210
rect 1920 -7260 2120 -7040
rect 1231 -7270 2120 -7260
rect 1231 -7340 1620 -7270
rect 1690 -7340 1930 -7270
rect 2000 -7340 2120 -7270
rect 1231 -7405 2120 -7340
rect 515 -7460 2120 -7405
rect 2290 -7295 2490 -6825
rect 2582 -6874 2636 -6864
rect 2582 -7028 2636 -7018
rect 2898 -6874 2952 -6864
rect 2898 -7028 2952 -7018
rect 3214 -6874 3268 -6864
rect 3214 -7028 3268 -7018
rect 2740 -7106 2794 -7096
rect 2740 -7260 2794 -7250
rect 3056 -7106 3110 -7096
rect 3056 -7260 3110 -7250
rect 3340 -7295 3540 -6825
rect 515 -7605 554 -7460
rect 754 -7540 1290 -7460
rect 1370 -7540 1431 -7460
rect 548 -7660 554 -7605
rect 754 -7605 1431 -7540
rect 754 -7660 760 -7605
rect 1914 -7660 1920 -7460
rect 2120 -7660 2126 -7460
rect 2290 -7500 3540 -7295
rect 4470 -6825 6142 -6620
rect 4470 -7295 4670 -6825
rect 4782 -6874 4836 -6864
rect 4782 -7028 4836 -7018
rect 5098 -6874 5152 -6864
rect 5098 -7028 5152 -7018
rect 5414 -6874 5468 -6864
rect 5414 -7028 5468 -7018
rect 4940 -7106 4994 -7096
rect 4940 -7260 4994 -7250
rect 5256 -7106 5310 -7096
rect 5256 -7260 5310 -7250
rect 5500 -7295 5700 -6825
rect 6350 -7290 7150 -20
rect 4470 -7500 5700 -7295
rect 1920 -7666 2120 -7660
rect 6344 -8090 6350 -7290
rect 7150 -8090 7156 -7290
rect 6350 -8096 7150 -8090
<< via1 >>
rect -270 2730 530 3530
rect 1630 2924 1830 2930
rect 1630 2736 1636 2924
rect 1636 2736 1824 2924
rect 1824 2736 1830 2924
rect 1630 2730 1830 2736
rect 2860 2730 3660 3530
rect 4650 2924 4850 2930
rect 4650 2736 4656 2924
rect 4656 2736 4844 2924
rect 4844 2736 4850 2924
rect 4650 2730 4850 2736
rect 6350 2730 7150 3530
rect 728 1727 933 1932
rect 2330 1730 2530 1930
rect 1940 940 2140 1140
rect 1110 580 1310 780
rect 2118 -1133 2323 -928
rect 3960 1730 4160 1930
rect 5510 1730 5710 1930
rect 4350 940 4550 1140
rect 4960 940 5160 1140
rect 4650 774 4850 780
rect 4650 586 4656 774
rect 4656 586 4844 774
rect 4844 586 4850 774
rect 4650 580 4850 586
rect 4350 -390 4550 -190
rect 4960 -740 5160 -540
rect 2860 -936 3660 -930
rect 2860 -1724 2866 -936
rect 2866 -1724 3654 -936
rect 3654 -1724 3660 -936
rect 3918 -1133 4123 -928
rect 2860 -1730 3660 -1724
rect 6350 -20 7150 780
rect 1192 -2319 1246 -2175
rect 1508 -2319 1562 -2175
rect 1824 -2319 1878 -2175
rect 1350 -2551 1404 -2407
rect 1666 -2551 1720 -2407
rect 2572 -2319 2626 -2175
rect 2888 -2319 2942 -2175
rect 3204 -2319 3258 -2175
rect 2730 -2551 2784 -2407
rect 3046 -2551 3100 -2407
rect 4742 -2319 4796 -2175
rect 5058 -2319 5112 -2175
rect 5374 -2319 5428 -2175
rect 4900 -2551 4954 -2407
rect 5216 -2551 5270 -2407
rect 5937 -1133 6142 -928
rect 2118 -6703 2323 -6498
rect 910 -7210 1030 -7090
rect 1750 -7210 1870 -7090
rect 2582 -7018 2636 -6874
rect 2898 -7018 2952 -6874
rect 3214 -7018 3268 -6874
rect 2740 -7250 2794 -7106
rect 3056 -7250 3110 -7106
rect 554 -7540 580 -7460
rect 580 -7540 660 -7460
rect 660 -7540 754 -7460
rect 554 -7660 754 -7540
rect 1920 -7466 2120 -7460
rect 1920 -7654 1926 -7466
rect 1926 -7654 2114 -7466
rect 2114 -7654 2120 -7466
rect 1920 -7660 2120 -7654
rect 4782 -7018 4836 -6874
rect 5098 -7018 5152 -6874
rect 5414 -7018 5468 -6874
rect 4940 -7250 4994 -7106
rect 5256 -7250 5310 -7106
rect 6350 -8090 7150 -7290
<< metal2 >>
rect 2860 3530 3660 3536
rect -470 2730 -270 3530
rect 530 2930 2860 3530
rect 530 2730 1630 2930
rect 1830 2730 2860 2930
rect 3660 2930 4860 3530
rect 3660 2730 4650 2930
rect 4850 2730 4860 2930
rect 6344 2730 6350 3530
rect 7150 2730 7156 3530
rect -270 2724 -70 2730
rect 1630 2500 1830 2730
rect 2860 2724 3660 2730
rect 4650 2500 4850 2730
rect 728 1932 933 1938
rect 933 1727 1172 1932
rect 2330 1930 2530 1936
rect 2250 1730 2330 1930
rect 728 1721 933 1727
rect 2330 1724 2530 1730
rect 3960 1930 4160 1936
rect 4160 1730 4240 1930
rect 5270 1730 5510 1930
rect 5710 1730 5716 1930
rect 3960 1724 4160 1730
rect 1940 1140 2140 1146
rect -470 940 1530 1140
rect 1110 780 1310 786
rect -470 580 1110 780
rect 1110 574 1310 580
rect 1630 780 1830 1120
rect 1940 934 2140 940
rect 4350 1140 4550 1146
rect 4960 1140 5160 1146
rect 4350 934 4550 940
rect 4650 780 4850 1140
rect 4960 934 5160 940
rect 6350 780 7150 786
rect 1630 580 4650 780
rect 4850 580 6350 780
rect 1630 -20 6350 580
rect 6350 -26 7150 -20
rect 4350 -190 4550 -184
rect -470 -390 4350 -190
rect 4350 -396 4550 -390
rect -470 -740 4960 -540
rect 5160 -740 5166 -540
rect 2118 -928 2323 -922
rect 3918 -928 4123 -922
rect -470 -2175 1890 -2130
rect -470 -2319 1192 -2175
rect 1246 -2319 1508 -2175
rect 1562 -2319 1824 -2175
rect 1878 -2319 1890 -2175
rect -470 -2330 1890 -2319
rect 1170 -2407 1890 -2400
rect 1170 -2530 1350 -2407
rect -470 -2551 1350 -2530
rect 1404 -2551 1666 -2407
rect 1720 -2551 1890 -2407
rect -470 -2600 1890 -2551
rect -470 -2730 1370 -2600
rect 2118 -6498 2323 -1133
rect 2854 -1530 2860 -930
rect 2560 -1730 2860 -1530
rect 3660 -1530 3666 -930
rect 4123 -1133 5937 -928
rect 6142 -1133 6148 -928
rect 3918 -1139 4123 -1133
rect 3660 -1730 5440 -1530
rect 2560 -2175 5440 -1730
rect 2560 -2319 2572 -2175
rect 2626 -2319 2888 -2175
rect 2942 -2319 3204 -2175
rect 3258 -2319 4742 -2175
rect 4796 -2319 5058 -2175
rect 5112 -2319 5374 -2175
rect 5428 -2319 5440 -2175
rect 2560 -2330 5440 -2319
rect 2560 -2407 3360 -2400
rect 2560 -2551 2730 -2407
rect 2784 -2551 3046 -2407
rect 3100 -2551 3360 -2407
rect 2560 -3660 3360 -2551
rect 4730 -2407 7950 -2400
rect 4730 -2551 4900 -2407
rect 4954 -2551 5216 -2407
rect 5270 -2551 7950 -2407
rect 4730 -3200 7950 -2551
rect 2560 -4460 7950 -3660
rect 2118 -6709 2323 -6703
rect 2570 -5740 7950 -4940
rect 2570 -6874 3370 -5740
rect 2570 -7018 2582 -6874
rect 2636 -7018 2898 -6874
rect 2952 -7018 3214 -6874
rect 3268 -7018 3370 -6874
rect 2570 -7030 3370 -7018
rect 4770 -6874 7950 -6230
rect 4770 -7018 4782 -6874
rect 4836 -7018 5098 -6874
rect 5152 -7018 5414 -6874
rect 5468 -7018 7950 -6874
rect 4770 -7030 7950 -7018
rect 871 -7050 1071 -7049
rect -470 -7090 1910 -7050
rect -470 -7210 910 -7090
rect 1030 -7210 1750 -7090
rect 1870 -7210 1910 -7090
rect -470 -7250 1910 -7210
rect 2570 -7106 5490 -7100
rect 2570 -7250 2740 -7106
rect 2794 -7250 3056 -7106
rect 3110 -7250 4940 -7106
rect 4994 -7250 5256 -7106
rect 5310 -7250 5490 -7106
rect 2570 -7290 5490 -7250
rect 6350 -7290 7150 -7284
rect 554 -7460 754 -7454
rect 1920 -7460 2120 -7454
rect 2570 -7460 6350 -7290
rect -470 -7660 554 -7460
rect 754 -7660 1920 -7460
rect 2120 -7660 6350 -7460
rect -470 -7900 6350 -7660
rect -470 -8260 3370 -7900
rect 4690 -8090 6350 -7900
rect 7150 -8090 7156 -7290
rect 6350 -8096 7150 -8090
use level_shifter_ad  level_shifter_ad_0
timestamp 1713664529
transform 1 0 140 0 1 2910
box 880 -1970 2310 -210
use level_shifter_ad  level_shifter_ad_1
timestamp 1713664529
transform 1 0 3160 0 1 2910
box 880 -1970 2310 -210
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_0
timestamp 1713663797
transform 1 0 973 0 1 -7147
box -423 -423 423 423
use sky130_fd_pr__diode_pw2nd_11v0_FT76RJ  sky130_fd_pr__diode_pw2nd_11v0_FT76RJ_0
timestamp 1713663180
transform 1 0 1812 0 1 -7147
box -217 -217 217 217
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM1
timestamp 1713252812
transform 1 0 5085 0 1 -2363
box -545 -497 545 497
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM2
timestamp 1713252812
transform 1 0 1535 0 1 -2363
box -545 -497 545 497
use sky130_fd_pr__nfet_g5v0d10v5_F7BQJ6  XM3
timestamp 1713252812
transform 1 0 5125 0 1 -7062
box -515 -458 515 458
use sky130_fd_pr__nfet_g5v0d10v5_F7BQJ6  XM21
timestamp 1713252812
transform 1 0 2925 0 1 -7062
box -515 -458 515 458
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM25
timestamp 1713252812
transform 1 0 2915 0 1 -2363
box -545 -497 545 497
<< labels >>
flabel metal2 -470 -2730 -270 -2530 0 FreeSans 256 0 0 0 EG_IBIAS
port 10 nsew
flabel metal2 -470 -2330 -270 -2130 0 FreeSans 256 0 0 0 IBIAS
port 5 nsew
flabel metal2 -470 -390 -270 -190 0 FreeSans 256 0 0 0 STDBY
port 4 nsew
flabel metal2 -470 -740 -270 -540 0 FreeSans 256 0 0 0 STDBY_B
port 13 nsew
flabel metal2 7150 -7030 7950 -6230 0 FreeSans 256 0 0 0 SG_AVSS
port 9 nsew
flabel metal2 7150 -5740 7950 -4940 0 FreeSans 256 0 0 0 EG_AVSS
port 7 nsew
flabel metal2 7150 -4460 7950 -3660 0 FreeSans 256 0 0 0 EG_AVDD
port 6 nsew
flabel metal2 7150 -3200 7950 -2400 0 FreeSans 256 0 0 0 SG_AVDD
port 8 nsew
flabel metal2 -470 -7250 -270 -7050 0 FreeSans 256 0 0 0 XIN
port 11 nsew
flabel metal2 -470 -8260 330 -7460 0 FreeSans 256 0 0 0 AVSS
port 2 nsew
flabel metal2 -470 580 -270 780 0 FreeSans 256 0 0 0 ENA_B
port 12 nsew
flabel metal2 -470 940 -270 1140 0 FreeSans 256 0 0 0 ENA
port 3 nsew
flabel metal2 -470 2730 330 3530 0 FreeSans 256 0 0 0 AVDD
port 1 nsew
flabel metal2 6350 2730 7150 3530 0 FreeSans 256 0 0 0 AVSS
port 2 nsew
<< end >>
