magic
tech sky130A
magscale 1 2
timestamp 1713441789
<< pwell >>
rect 1560 -1860 1630 -1144
<< locali >>
rect 1044 -360 1532 -354
rect 1654 -360 2142 -354
rect 1038 -428 1538 -360
rect 1038 -958 1112 -428
rect 1464 -470 1538 -428
rect 1464 -916 1484 -470
rect 1518 -916 1538 -470
rect 1464 -958 1538 -916
rect 1038 -1026 1538 -958
rect 1648 -428 2148 -360
rect 1648 -470 1722 -428
rect 1648 -916 1668 -470
rect 1702 -916 1722 -470
rect 1648 -958 1722 -916
rect 2074 -958 2148 -428
rect 1648 -1026 2148 -958
rect 1044 -1032 1532 -1026
rect 1654 -1032 2142 -1026
rect 1044 -1178 1532 -1172
rect 1654 -1178 2142 -1172
rect 1038 -1246 1538 -1178
rect 1038 -1758 1112 -1246
rect 1464 -1288 1538 -1246
rect 1464 -1716 1484 -1288
rect 1518 -1716 1538 -1288
rect 1464 -1758 1538 -1716
rect 1038 -1826 1538 -1758
rect 1648 -1246 2148 -1178
rect 1648 -1288 1722 -1246
rect 1648 -1716 1668 -1288
rect 1702 -1716 1722 -1288
rect 1648 -1758 1722 -1716
rect 2074 -1758 2148 -1246
rect 1648 -1826 2148 -1758
rect 1044 -1832 1532 -1826
rect 1654 -1832 2142 -1826
<< viali >>
rect 1484 -916 1518 -470
rect 1668 -916 1702 -470
rect 1484 -1716 1518 -1288
rect 1668 -1716 1702 -1288
<< metal1 >>
rect 1540 -260 1640 -254
rect 1540 -450 1640 -360
rect 1232 -560 1238 -460
rect 1338 -560 1344 -460
rect 1464 -470 1722 -450
rect 1464 -643 1484 -470
rect 1030 -743 1226 -643
rect 1350 -743 1484 -643
rect 1030 -1030 1130 -743
rect 1232 -930 1238 -830
rect 1338 -930 1344 -830
rect 1464 -916 1484 -743
rect 1518 -743 1668 -470
rect 1518 -916 1538 -743
rect 1464 -936 1538 -916
rect 1648 -916 1668 -743
rect 1702 -643 1722 -470
rect 1842 -560 1848 -460
rect 1948 -560 1954 -460
rect 1702 -743 1836 -643
rect 1954 -743 2160 -643
rect 1702 -916 1722 -743
rect 1648 -936 1722 -916
rect 1848 -830 1948 -824
rect 1948 -930 1954 -830
rect 1848 -1030 1948 -930
rect 1024 -1130 1030 -1030
rect 1130 -1130 1948 -1030
rect 2060 -1030 2160 -743
rect 1030 -1452 1130 -1130
rect 1232 -1370 1238 -1270
rect 1338 -1370 1344 -1270
rect 1464 -1288 1538 -1268
rect 1464 -1452 1484 -1288
rect 1030 -1552 1226 -1452
rect 1350 -1552 1484 -1452
rect 1232 -1730 1238 -1630
rect 1338 -1730 1344 -1630
rect 1464 -1716 1484 -1552
rect 1518 -1452 1538 -1288
rect 1648 -1288 1722 -1268
rect 1648 -1452 1668 -1288
rect 1518 -1716 1668 -1452
rect 1702 -1452 1722 -1288
rect 1842 -1370 1848 -1270
rect 1948 -1370 1954 -1270
rect 2060 -1452 2160 -1130
rect 1702 -1552 1836 -1452
rect 1954 -1552 2160 -1452
rect 1702 -1716 1722 -1552
rect 1464 -1736 1722 -1716
rect 1844 -1730 1850 -1630
rect 1950 -1730 1956 -1630
rect 1540 -1820 1640 -1736
rect 1540 -1926 1640 -1920
<< via1 >>
rect 1540 -360 1640 -260
rect 1238 -560 1338 -460
rect 1238 -930 1338 -830
rect 1848 -560 1948 -460
rect 1848 -930 1948 -830
rect 1030 -1130 1130 -1030
rect 2060 -1130 2160 -1030
rect 1238 -1370 1338 -1270
rect 1238 -1730 1338 -1630
rect 1848 -1370 1948 -1270
rect 1850 -1730 1950 -1630
rect 1540 -1920 1640 -1820
<< metal2 >>
rect 1490 -260 1690 -210
rect 1490 -360 1540 -260
rect 1640 -360 1690 -260
rect 1490 -410 1690 -360
rect 1238 -460 1338 -454
rect 1238 -830 1338 -560
rect 1848 -460 1948 -454
rect 1848 -830 1948 -560
rect 1338 -930 1340 -830
rect 1842 -930 1848 -830
rect 1948 -930 1954 -830
rect 880 -1024 1080 -980
rect 880 -1030 1130 -1024
rect 880 -1130 1030 -1030
rect 1238 -1030 1338 -930
rect 1848 -936 1948 -930
rect 2110 -1030 2310 -980
rect 1238 -1130 2060 -1030
rect 2160 -1130 2310 -1030
rect 880 -1136 1130 -1130
rect 880 -1180 1080 -1136
rect 2110 -1180 2310 -1130
rect 1238 -1270 1338 -1264
rect 1238 -1630 1338 -1370
rect 1238 -1770 1338 -1730
rect 1848 -1270 1948 -1264
rect 1948 -1370 1950 -1297
rect 1848 -1630 1950 -1370
rect 1848 -1730 1850 -1630
rect 1848 -1770 1950 -1730
rect 1190 -1970 1390 -1770
rect 1490 -1820 1690 -1770
rect 1490 -1920 1540 -1820
rect 1640 -1920 1690 -1820
rect 1490 -1970 1690 -1920
rect 1800 -1970 2000 -1770
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM1
timestamp 1713252812
transform 1 0 1898 0 1 -693
box -308 -397 308 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM2
timestamp 1713441789
transform 1 0 1898 0 1 -1502
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM21
timestamp 1713441789
transform 1 0 1288 0 1 -1502
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM25
timestamp 1713252812
transform 1 0 1288 0 1 -693
box -308 -397 308 397
<< labels >>
flabel metal2 1490 -410 1690 -210 0 FreeSans 256 0 0 0 AVDD
port 1 nsew
flabel metal2 880 -1180 1080 -980 0 FreeSans 256 0 0 0 HI_B
port 5 nsew
flabel metal2 1190 -1970 1390 -1770 0 FreeSans 256 0 0 0 LO
port 2 nsew
flabel metal2 1800 -1970 2000 -1770 0 FreeSans 256 0 0 0 LO_B
port 3 nsew
flabel metal2 1490 -1970 1690 -1770 0 FreeSans 256 0 0 0 AVSS
port 0 nsew
flabel metal2 2110 -1180 2310 -980 0 FreeSans 256 0 0 0 HI
port 4 nsew
<< end >>
