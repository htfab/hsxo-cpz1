magic
tech sky130A
magscale 1 2
timestamp 1713747467
<< nwell >>
rect -545 -3497 545 3497
<< mvpmos >>
rect -287 -3200 -187 3200
rect -129 -3200 -29 3200
rect 29 -3200 129 3200
rect 187 -3200 287 3200
<< mvpdiff >>
rect -345 3188 -287 3200
rect -345 -3188 -333 3188
rect -299 -3188 -287 3188
rect -345 -3200 -287 -3188
rect -187 3188 -129 3200
rect -187 -3188 -175 3188
rect -141 -3188 -129 3188
rect -187 -3200 -129 -3188
rect -29 3188 29 3200
rect -29 -3188 -17 3188
rect 17 -3188 29 3188
rect -29 -3200 29 -3188
rect 129 3188 187 3200
rect 129 -3188 141 3188
rect 175 -3188 187 3188
rect 129 -3200 187 -3188
rect 287 3188 345 3200
rect 287 -3188 299 3188
rect 333 -3188 345 3188
rect 287 -3200 345 -3188
<< mvpdiffc >>
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
<< mvnsubdiff >>
rect -479 3419 479 3431
rect -479 3385 -371 3419
rect 371 3385 479 3419
rect -479 3373 479 3385
rect -479 3323 -421 3373
rect -479 -3323 -467 3323
rect -433 -3323 -421 3323
rect 421 3323 479 3373
rect -479 -3373 -421 -3323
rect 421 -3323 433 3323
rect 467 -3323 479 3323
rect 421 -3373 479 -3323
rect -479 -3385 479 -3373
rect -479 -3419 -371 -3385
rect 371 -3419 479 -3385
rect -479 -3431 479 -3419
<< mvnsubdiffcont >>
rect -371 3385 371 3419
rect -467 -3323 -433 3323
rect 433 -3323 467 3323
rect -371 -3419 371 -3385
<< poly >>
rect -287 3281 -187 3297
rect -287 3247 -271 3281
rect -203 3247 -187 3281
rect -287 3200 -187 3247
rect -129 3281 -29 3297
rect -129 3247 -113 3281
rect -45 3247 -29 3281
rect -129 3200 -29 3247
rect 29 3281 129 3297
rect 29 3247 45 3281
rect 113 3247 129 3281
rect 29 3200 129 3247
rect 187 3281 287 3297
rect 187 3247 203 3281
rect 271 3247 287 3281
rect 187 3200 287 3247
rect -287 -3247 -187 -3200
rect -287 -3281 -271 -3247
rect -203 -3281 -187 -3247
rect -287 -3297 -187 -3281
rect -129 -3247 -29 -3200
rect -129 -3281 -113 -3247
rect -45 -3281 -29 -3247
rect -129 -3297 -29 -3281
rect 29 -3247 129 -3200
rect 29 -3281 45 -3247
rect 113 -3281 129 -3247
rect 29 -3297 129 -3281
rect 187 -3247 287 -3200
rect 187 -3281 203 -3247
rect 271 -3281 287 -3247
rect 187 -3297 287 -3281
<< polycont >>
rect -271 3247 -203 3281
rect -113 3247 -45 3281
rect 45 3247 113 3281
rect 203 3247 271 3281
rect -271 -3281 -203 -3247
rect -113 -3281 -45 -3247
rect 45 -3281 113 -3247
rect 203 -3281 271 -3247
<< locali >>
rect -467 3385 -371 3419
rect 371 3385 467 3419
rect -467 3323 -433 3385
rect 433 3323 467 3385
rect -287 3247 -271 3281
rect -203 3247 -187 3281
rect -129 3247 -113 3281
rect -45 3247 -29 3281
rect 29 3247 45 3281
rect 113 3247 129 3281
rect 187 3247 203 3281
rect 271 3247 287 3281
rect -333 3188 -299 3204
rect -333 -3204 -299 -3188
rect -175 3188 -141 3204
rect -175 -3204 -141 -3188
rect -17 3188 17 3204
rect -17 -3204 17 -3188
rect 141 3188 175 3204
rect 141 -3204 175 -3188
rect 299 3188 333 3204
rect 299 -3204 333 -3188
rect -287 -3281 -271 -3247
rect -203 -3281 -187 -3247
rect -129 -3281 -113 -3247
rect -45 -3281 -29 -3247
rect 29 -3281 45 -3247
rect 113 -3281 129 -3247
rect 187 -3281 203 -3247
rect 271 -3281 287 -3247
rect -467 -3385 -433 -3323
rect 433 -3385 467 -3323
rect -467 -3419 -371 -3385
rect 371 -3419 467 -3385
<< viali >>
rect -271 3247 -203 3281
rect -113 3247 -45 3281
rect 45 3247 113 3281
rect 203 3247 271 3281
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
rect -271 -3281 -203 -3247
rect -113 -3281 -45 -3247
rect 45 -3281 113 -3247
rect 203 -3281 271 -3247
<< metal1 >>
rect -283 3281 -191 3287
rect -283 3247 -271 3281
rect -203 3247 -191 3281
rect -283 3241 -191 3247
rect -125 3281 -33 3287
rect -125 3247 -113 3281
rect -45 3247 -33 3281
rect -125 3241 -33 3247
rect 33 3281 125 3287
rect 33 3247 45 3281
rect 113 3247 125 3281
rect 33 3241 125 3247
rect 191 3281 283 3287
rect 191 3247 203 3281
rect 271 3247 283 3281
rect 191 3241 283 3247
rect -339 3188 -293 3200
rect -339 -3188 -333 3188
rect -299 -3188 -293 3188
rect -339 -3200 -293 -3188
rect -181 3188 -135 3200
rect -181 -3188 -175 3188
rect -141 -3188 -135 3188
rect -181 -3200 -135 -3188
rect -23 3188 23 3200
rect -23 -3188 -17 3188
rect 17 -3188 23 3188
rect -23 -3200 23 -3188
rect 135 3188 181 3200
rect 135 -3188 141 3188
rect 175 -3188 181 3188
rect 135 -3200 181 -3188
rect 293 3188 339 3200
rect 293 -3188 299 3188
rect 333 -3188 339 3188
rect 293 -3200 339 -3188
rect -283 -3247 -191 -3241
rect -283 -3281 -271 -3247
rect -203 -3281 -191 -3247
rect -283 -3287 -191 -3281
rect -125 -3247 -33 -3241
rect -125 -3281 -113 -3247
rect -45 -3281 -33 -3247
rect -125 -3287 -33 -3281
rect 33 -3247 125 -3241
rect 33 -3281 45 -3247
rect 113 -3281 125 -3247
rect 33 -3287 125 -3281
rect 191 -3247 283 -3241
rect 191 -3281 203 -3247
rect 271 -3281 283 -3247
rect 191 -3287 283 -3281
<< properties >>
string FIXED_BBOX -450 -3402 450 3402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
