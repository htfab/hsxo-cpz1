magic
tech sky130A
magscale 1 2
timestamp 1712784051
<< pwell >>
rect -201 -2182 201 2182
<< psubdiff >>
rect -165 2112 -69 2146
rect 69 2112 165 2146
rect -165 2050 -131 2112
rect 131 2050 165 2112
rect -165 -2112 -131 -2050
rect 131 -2112 165 -2050
rect -165 -2146 -69 -2112
rect 69 -2146 165 -2112
<< psubdiffcont >>
rect -69 2112 69 2146
rect -165 -2050 -131 2050
rect 131 -2050 165 2050
rect -69 -2146 69 -2112
<< xpolycontact >>
rect -35 1584 35 2016
rect -35 -2016 35 -1584
<< xpolyres >>
rect -35 -1584 35 1584
<< locali >>
rect -165 2112 -69 2146
rect 69 2112 165 2146
rect -165 2050 -131 2112
rect 131 2050 165 2112
rect -165 -2112 -131 -2050
rect 131 -2112 165 -2050
rect -165 -2146 -69 -2112
rect 69 -2146 165 -2112
<< viali >>
rect -19 1601 19 1998
rect -19 -1998 19 -1601
<< metal1 >>
rect -25 1998 25 2010
rect -25 1601 -19 1998
rect 19 1601 25 1998
rect -25 1589 25 1601
rect -25 -1601 25 -1589
rect -25 -1998 -19 -1601
rect 19 -1998 25 -1601
rect -25 -2010 25 -1998
<< properties >>
string FIXED_BBOX -148 -2129 148 2129
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 16.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 92.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
