magic
tech sky130A
magscale 1 2
timestamp 1713804741
<< error_p >>
rect -269 472 -211 478
rect -77 472 -19 478
rect 115 472 173 478
rect 307 472 365 478
rect -269 438 -257 472
rect -77 438 -65 472
rect 115 438 127 472
rect 307 438 319 472
rect -269 432 -211 438
rect -77 432 -19 438
rect 115 432 173 438
rect 307 432 365 438
rect -365 -438 -307 -432
rect -173 -438 -115 -432
rect 19 -438 77 -432
rect 211 -438 269 -432
rect -365 -472 -353 -438
rect -173 -472 -161 -438
rect 19 -472 31 -438
rect 211 -472 223 -438
rect -365 -478 -307 -472
rect -173 -478 -115 -472
rect 19 -478 77 -472
rect 211 -478 269 -472
<< pwell >>
rect -551 -610 551 610
<< nmos >>
rect -351 -400 -321 400
rect -255 -400 -225 400
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
rect 225 -400 255 400
rect 321 -400 351 400
<< ndiff >>
rect -413 388 -351 400
rect -413 -388 -401 388
rect -367 -388 -351 388
rect -413 -400 -351 -388
rect -321 388 -255 400
rect -321 -388 -305 388
rect -271 -388 -255 388
rect -321 -400 -255 -388
rect -225 388 -159 400
rect -225 -388 -209 388
rect -175 -388 -159 388
rect -225 -400 -159 -388
rect -129 388 -63 400
rect -129 -388 -113 388
rect -79 -388 -63 388
rect -129 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 129 400
rect 63 -388 79 388
rect 113 -388 129 388
rect 63 -400 129 -388
rect 159 388 225 400
rect 159 -388 175 388
rect 209 -388 225 388
rect 159 -400 225 -388
rect 255 388 321 400
rect 255 -388 271 388
rect 305 -388 321 388
rect 255 -400 321 -388
rect 351 388 413 400
rect 351 -388 367 388
rect 401 -388 413 388
rect 351 -400 413 -388
<< ndiffc >>
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
<< psubdiff >>
rect -515 540 -419 574
rect 419 540 515 574
rect -515 478 -481 540
rect 481 478 515 540
rect -515 -540 -481 -478
rect 481 -540 515 -478
rect -515 -574 -419 -540
rect 419 -574 515 -540
<< psubdiffcont >>
rect -419 540 419 574
rect -515 -478 -481 478
rect 481 -478 515 478
rect -419 -574 419 -540
<< poly >>
rect -273 472 -207 488
rect -273 438 -257 472
rect -223 438 -207 472
rect -351 400 -321 426
rect -273 422 -207 438
rect -81 472 -15 488
rect -81 438 -65 472
rect -31 438 -15 472
rect -255 400 -225 422
rect -159 400 -129 426
rect -81 422 -15 438
rect 111 472 177 488
rect 111 438 127 472
rect 161 438 177 472
rect -63 400 -33 422
rect 33 400 63 426
rect 111 422 177 438
rect 303 472 369 488
rect 303 438 319 472
rect 353 438 369 472
rect 129 400 159 422
rect 225 400 255 426
rect 303 422 369 438
rect 321 400 351 422
rect -351 -422 -321 -400
rect -369 -438 -303 -422
rect -255 -426 -225 -400
rect -159 -422 -129 -400
rect -369 -472 -353 -438
rect -319 -472 -303 -438
rect -369 -488 -303 -472
rect -177 -438 -111 -422
rect -63 -426 -33 -400
rect 33 -422 63 -400
rect -177 -472 -161 -438
rect -127 -472 -111 -438
rect -177 -488 -111 -472
rect 15 -438 81 -422
rect 129 -426 159 -400
rect 225 -422 255 -400
rect 15 -472 31 -438
rect 65 -472 81 -438
rect 15 -488 81 -472
rect 207 -438 273 -422
rect 321 -426 351 -400
rect 207 -472 223 -438
rect 257 -472 273 -438
rect 207 -488 273 -472
<< polycont >>
rect -257 438 -223 472
rect -65 438 -31 472
rect 127 438 161 472
rect 319 438 353 472
rect -353 -472 -319 -438
rect -161 -472 -127 -438
rect 31 -472 65 -438
rect 223 -472 257 -438
<< locali >>
rect -515 540 -419 574
rect 419 540 515 574
rect -515 478 -481 540
rect 481 478 515 540
rect -273 438 -257 472
rect -223 438 -207 472
rect -81 438 -65 472
rect -31 438 -15 472
rect 111 438 127 472
rect 161 438 177 472
rect 303 438 319 472
rect 353 438 369 472
rect -401 388 -367 404
rect -401 -404 -367 -388
rect -305 388 -271 404
rect -305 -404 -271 -388
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect 271 388 305 404
rect 271 -404 305 -388
rect 367 388 401 404
rect 367 -404 401 -388
rect -369 -472 -353 -438
rect -319 -472 -303 -438
rect -177 -472 -161 -438
rect -127 -472 -111 -438
rect 15 -472 31 -438
rect 65 -472 81 -438
rect 207 -472 223 -438
rect 257 -472 273 -438
rect -515 -540 -481 -478
rect 481 -540 515 -478
rect -515 -574 -419 -540
rect 419 -574 515 -540
<< viali >>
rect -257 438 -223 472
rect -65 438 -31 472
rect 127 438 161 472
rect 319 438 353 472
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
rect -353 -472 -319 -438
rect -161 -472 -127 -438
rect 31 -472 65 -438
rect 223 -472 257 -438
<< metal1 >>
rect -269 472 -211 478
rect -269 438 -257 472
rect -223 438 -211 472
rect -269 432 -211 438
rect -77 472 -19 478
rect -77 438 -65 472
rect -31 438 -19 472
rect -77 432 -19 438
rect 115 472 173 478
rect 115 438 127 472
rect 161 438 173 472
rect 115 432 173 438
rect 307 472 365 478
rect 307 438 319 472
rect 353 438 365 472
rect 307 432 365 438
rect -407 388 -361 400
rect -407 -388 -401 388
rect -367 -388 -361 388
rect -407 -400 -361 -388
rect -311 388 -265 400
rect -311 -388 -305 388
rect -271 -388 -265 388
rect -311 -400 -265 -388
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect 265 388 311 400
rect 265 -388 271 388
rect 305 -388 311 388
rect 265 -400 311 -388
rect 361 388 407 400
rect 361 -388 367 388
rect 401 -388 407 388
rect 361 -400 407 -388
rect -365 -438 -307 -432
rect -365 -472 -353 -438
rect -319 -472 -307 -438
rect -365 -478 -307 -472
rect -173 -438 -115 -432
rect -173 -472 -161 -438
rect -127 -472 -115 -438
rect -173 -478 -115 -472
rect 19 -438 77 -432
rect 19 -472 31 -438
rect 65 -472 77 -438
rect 19 -478 77 -472
rect 211 -438 269 -432
rect 211 -472 223 -438
rect 257 -472 269 -438
rect 211 -478 269 -472
<< properties >>
string FIXED_BBOX -498 -557 498 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
