magic
tech sky130A
magscale 1 2
timestamp 1713747467
<< pwell >>
rect -515 -3458 515 3458
<< mvnmos >>
rect -287 -3200 -187 3200
rect -129 -3200 -29 3200
rect 29 -3200 129 3200
rect 187 -3200 287 3200
<< mvndiff >>
rect -345 3188 -287 3200
rect -345 -3188 -333 3188
rect -299 -3188 -287 3188
rect -345 -3200 -287 -3188
rect -187 3188 -129 3200
rect -187 -3188 -175 3188
rect -141 -3188 -129 3188
rect -187 -3200 -129 -3188
rect -29 3188 29 3200
rect -29 -3188 -17 3188
rect 17 -3188 29 3188
rect -29 -3200 29 -3188
rect 129 3188 187 3200
rect 129 -3188 141 3188
rect 175 -3188 187 3188
rect 129 -3200 187 -3188
rect 287 3188 345 3200
rect 287 -3188 299 3188
rect 333 -3188 345 3188
rect 287 -3200 345 -3188
<< mvndiffc >>
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
<< mvpsubdiff >>
rect -479 3410 479 3422
rect -479 3376 -371 3410
rect 371 3376 479 3410
rect -479 3364 479 3376
rect -479 3314 -421 3364
rect -479 -3314 -467 3314
rect -433 -3314 -421 3314
rect 421 3314 479 3364
rect -479 -3364 -421 -3314
rect 421 -3314 433 3314
rect 467 -3314 479 3314
rect 421 -3364 479 -3314
rect -479 -3376 479 -3364
rect -479 -3410 -371 -3376
rect 371 -3410 479 -3376
rect -479 -3422 479 -3410
<< mvpsubdiffcont >>
rect -371 3376 371 3410
rect -467 -3314 -433 3314
rect 433 -3314 467 3314
rect -371 -3410 371 -3376
<< poly >>
rect -287 3272 -187 3288
rect -287 3238 -271 3272
rect -203 3238 -187 3272
rect -287 3200 -187 3238
rect -129 3272 -29 3288
rect -129 3238 -113 3272
rect -45 3238 -29 3272
rect -129 3200 -29 3238
rect 29 3272 129 3288
rect 29 3238 45 3272
rect 113 3238 129 3272
rect 29 3200 129 3238
rect 187 3272 287 3288
rect 187 3238 203 3272
rect 271 3238 287 3272
rect 187 3200 287 3238
rect -287 -3238 -187 -3200
rect -287 -3272 -271 -3238
rect -203 -3272 -187 -3238
rect -287 -3288 -187 -3272
rect -129 -3238 -29 -3200
rect -129 -3272 -113 -3238
rect -45 -3272 -29 -3238
rect -129 -3288 -29 -3272
rect 29 -3238 129 -3200
rect 29 -3272 45 -3238
rect 113 -3272 129 -3238
rect 29 -3288 129 -3272
rect 187 -3238 287 -3200
rect 187 -3272 203 -3238
rect 271 -3272 287 -3238
rect 187 -3288 287 -3272
<< polycont >>
rect -271 3238 -203 3272
rect -113 3238 -45 3272
rect 45 3238 113 3272
rect 203 3238 271 3272
rect -271 -3272 -203 -3238
rect -113 -3272 -45 -3238
rect 45 -3272 113 -3238
rect 203 -3272 271 -3238
<< locali >>
rect -467 3376 -371 3410
rect 371 3376 467 3410
rect -467 3314 -433 3376
rect 433 3314 467 3376
rect -287 3238 -271 3272
rect -203 3238 -187 3272
rect -129 3238 -113 3272
rect -45 3238 -29 3272
rect 29 3238 45 3272
rect 113 3238 129 3272
rect 187 3238 203 3272
rect 271 3238 287 3272
rect -333 3188 -299 3204
rect -333 -3204 -299 -3188
rect -175 3188 -141 3204
rect -175 -3204 -141 -3188
rect -17 3188 17 3204
rect -17 -3204 17 -3188
rect 141 3188 175 3204
rect 141 -3204 175 -3188
rect 299 3188 333 3204
rect 299 -3204 333 -3188
rect -287 -3272 -271 -3238
rect -203 -3272 -187 -3238
rect -129 -3272 -113 -3238
rect -45 -3272 -29 -3238
rect 29 -3272 45 -3238
rect 113 -3272 129 -3238
rect 187 -3272 203 -3238
rect 271 -3272 287 -3238
rect -467 -3376 -433 -3314
rect 433 -3376 467 -3314
rect -467 -3410 -371 -3376
rect 371 -3410 467 -3376
<< viali >>
rect -271 3238 -203 3272
rect -113 3238 -45 3272
rect 45 3238 113 3272
rect 203 3238 271 3272
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
rect -271 -3272 -203 -3238
rect -113 -3272 -45 -3238
rect 45 -3272 113 -3238
rect 203 -3272 271 -3238
<< metal1 >>
rect -283 3272 -191 3278
rect -283 3238 -271 3272
rect -203 3238 -191 3272
rect -283 3232 -191 3238
rect -125 3272 -33 3278
rect -125 3238 -113 3272
rect -45 3238 -33 3272
rect -125 3232 -33 3238
rect 33 3272 125 3278
rect 33 3238 45 3272
rect 113 3238 125 3272
rect 33 3232 125 3238
rect 191 3272 283 3278
rect 191 3238 203 3272
rect 271 3238 283 3272
rect 191 3232 283 3238
rect -339 3188 -293 3200
rect -339 -3188 -333 3188
rect -299 -3188 -293 3188
rect -339 -3200 -293 -3188
rect -181 3188 -135 3200
rect -181 -3188 -175 3188
rect -141 -3188 -135 3188
rect -181 -3200 -135 -3188
rect -23 3188 23 3200
rect -23 -3188 -17 3188
rect 17 -3188 23 3188
rect -23 -3200 23 -3188
rect 135 3188 181 3200
rect 135 -3188 141 3188
rect 175 -3188 181 3188
rect 135 -3200 181 -3188
rect 293 3188 339 3200
rect 293 -3188 299 3188
rect 333 -3188 339 3188
rect 293 -3200 339 -3188
rect -283 -3238 -191 -3232
rect -283 -3272 -271 -3238
rect -203 -3272 -191 -3238
rect -283 -3278 -191 -3272
rect -125 -3238 -33 -3232
rect -125 -3272 -113 -3238
rect -45 -3272 -33 -3238
rect -125 -3278 -33 -3272
rect 33 -3238 125 -3232
rect 33 -3272 45 -3238
rect 113 -3272 125 -3238
rect 33 -3278 125 -3272
rect 191 -3238 283 -3232
rect 191 -3272 203 -3238
rect 271 -3272 283 -3238
rect 191 -3278 283 -3272
<< properties >>
string FIXED_BBOX -450 -3393 450 3393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
