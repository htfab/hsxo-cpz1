magic
tech sky130A
magscale 1 2
timestamp 1713792225
<< nwell >>
rect 1400 -3210 2070 -1720
rect 2490 -2360 4124 -1720
rect 1400 -4440 2100 -3210
<< pwell >>
rect 2500 -2980 4124 -2360
rect 3854 -4620 4544 -2980
rect 3854 -4710 4928 -4620
rect 3204 -5930 3854 -4710
<< locali >>
rect 2092 -1744 2470 -1738
rect 4146 -1744 4524 -1738
rect 2086 -1812 2476 -1744
rect 2086 -1940 2160 -1812
rect 1310 -2140 2160 -1940
rect 2086 -2270 2160 -2140
rect 2402 -2270 2476 -1812
rect 4140 -1812 4530 -1744
rect 4140 -1940 4214 -1812
rect 3584 -1946 4214 -1940
rect 3584 -2134 3590 -1946
rect 3778 -2134 4214 -1946
rect 3584 -2140 4214 -2134
rect 2086 -2338 2476 -2270
rect 4140 -2270 4214 -2140
rect 4456 -2270 4530 -1812
rect 4140 -2338 4530 -2270
rect 2092 -2340 2470 -2338
rect 4146 -2340 4524 -2338
rect 2092 -2382 2470 -2380
rect 4146 -2382 4524 -2380
rect 2086 -2450 2476 -2382
rect 2086 -2890 2160 -2450
rect 2402 -2890 2476 -2450
rect 4140 -2450 4530 -2382
rect 4140 -2760 4214 -2450
rect 2086 -2958 2476 -2890
rect 3964 -2890 4214 -2760
rect 4456 -2890 4530 -2450
rect 3964 -2958 4530 -2890
rect 2092 -2964 2470 -2958
rect 3964 -2964 4524 -2958
rect 3964 -3026 4164 -2964
rect 3964 -3214 3970 -3026
rect 4158 -3214 4164 -3026
rect 3964 -3220 4164 -3214
rect 2122 -3234 3180 -3228
rect 2116 -3302 3186 -3234
rect 2116 -3390 2190 -3302
rect 1510 -3396 2190 -3390
rect 1694 -3584 2190 -3396
rect 1510 -3590 2190 -3584
rect 2116 -4360 2190 -3590
rect 3112 -4360 3186 -3302
rect 2116 -4428 3186 -4360
rect 2122 -4434 3180 -4428
rect 2124 -4732 3182 -4726
rect 3876 -4732 4934 -4726
rect 2118 -4800 3188 -4732
rect 2118 -5840 2192 -4800
rect 3114 -5560 3188 -4800
rect 3870 -4800 4940 -4732
rect 3870 -5560 3944 -4800
rect 3114 -5760 3944 -5560
rect 3114 -5840 3188 -5760
rect 2118 -5908 3188 -5840
rect 3870 -5840 3944 -5760
rect 4866 -5560 4940 -4800
rect 4866 -5566 5558 -5560
rect 4866 -5754 5364 -5566
rect 5552 -5754 5558 -5566
rect 4866 -5760 5558 -5754
rect 4866 -5840 4940 -5760
rect 3870 -5908 4940 -5840
rect 2124 -5914 3182 -5908
rect 3876 -5914 4934 -5908
<< viali >>
rect 1110 -2140 1310 -1940
rect 3590 -2134 3778 -1946
rect 3970 -3214 4158 -3026
rect 1506 -3584 1694 -3396
rect 5364 -5754 5552 -5566
<< metal1 >>
rect 1494 -1720 1500 -1520
rect 1700 -1720 1706 -1520
rect 1104 -1940 1316 -1928
rect 1104 -2140 1110 -1940
rect 1310 -2140 1316 -1940
rect 1104 -2152 1316 -2140
rect 1110 -3390 1310 -2152
rect 1500 -2880 1700 -1720
rect 3584 -1940 3784 -1934
rect 3578 -2140 3584 -1940
rect 3784 -2140 3790 -1940
rect 3188 -2460 3194 -2260
rect 3394 -2460 3400 -2260
rect 1494 -3080 1500 -2880
rect 1700 -3080 1706 -2880
rect 3194 -3190 3394 -2460
rect 1500 -3390 1700 -3384
rect 1104 -3590 1110 -3390
rect 1310 -3590 1316 -3390
rect 1500 -3596 1700 -3590
rect 1900 -3390 3394 -3190
rect 1900 -4270 2100 -3390
rect 2240 -3443 2294 -3433
rect 2240 -3597 2294 -3587
rect 2432 -3443 2486 -3433
rect 2432 -3597 2486 -3587
rect 2624 -3443 2678 -3433
rect 2624 -3597 2678 -3587
rect 2816 -3443 2870 -3433
rect 2816 -3597 2870 -3587
rect 3008 -3443 3062 -3433
rect 3008 -3597 3062 -3587
rect 2336 -4075 2390 -4065
rect 2336 -4229 2390 -4219
rect 2528 -4075 2582 -4065
rect 2528 -4229 2582 -4219
rect 2720 -4075 2774 -4065
rect 2720 -4229 2774 -4219
rect 2912 -4075 2966 -4065
rect 2912 -4229 2966 -4219
rect 3194 -4270 3394 -3390
rect 3584 -3390 3784 -2140
rect 4704 -2260 4904 -2254
rect 3958 -3220 3964 -3020
rect 4164 -3220 4170 -3020
rect 4704 -3040 4904 -2460
rect 3584 -3596 3784 -3590
rect 4504 -3240 4904 -3040
rect 1500 -4470 3854 -4270
rect 1500 -4490 1700 -4470
rect 3196 -4690 3396 -4684
rect 1500 -4696 1700 -4690
rect 1902 -4890 3196 -4690
rect 1902 -5760 2102 -4890
rect 2242 -4932 2296 -4922
rect 2242 -5086 2296 -5076
rect 2434 -4932 2488 -4922
rect 2434 -5086 2488 -5076
rect 2626 -4932 2680 -4922
rect 2626 -5086 2680 -5076
rect 2818 -4932 2872 -4922
rect 2818 -5086 2872 -5076
rect 3010 -4932 3064 -4922
rect 3010 -5086 3064 -5076
rect 2338 -5564 2392 -5554
rect 2338 -5718 2392 -5708
rect 2530 -5564 2584 -5554
rect 2530 -5718 2584 -5708
rect 2722 -5564 2776 -5554
rect 2722 -5718 2776 -5708
rect 2914 -5564 2968 -5554
rect 2914 -5718 2968 -5708
rect 3196 -5760 3396 -4890
rect 1500 -5960 3396 -5760
rect 3654 -4690 3854 -4470
rect 4504 -4370 4704 -3240
rect 5352 -3660 5358 -3460
rect 5558 -3660 5564 -3460
rect 4504 -4576 4704 -4570
rect 3654 -4890 5158 -4690
rect 3654 -5750 3854 -4890
rect 3994 -4932 4048 -4922
rect 3994 -5086 4048 -5076
rect 4186 -4932 4240 -4922
rect 4186 -5086 4240 -5076
rect 4378 -4932 4432 -4922
rect 4378 -5086 4432 -5076
rect 4570 -4932 4624 -4922
rect 4570 -5086 4624 -5076
rect 4762 -4932 4816 -4922
rect 4762 -5086 4816 -5076
rect 4090 -5564 4144 -5554
rect 4090 -5718 4144 -5708
rect 4282 -5564 4336 -5554
rect 4282 -5718 4336 -5708
rect 4474 -5564 4528 -5554
rect 4474 -5718 4528 -5708
rect 4666 -5564 4720 -5554
rect 4666 -5718 4720 -5708
rect 4958 -5750 5158 -4890
rect 3654 -5960 5158 -5750
rect 5358 -5560 5558 -3660
rect 5358 -5766 5558 -5760
rect 1500 -5980 1700 -5960
rect 1500 -6186 1700 -6180
<< via1 >>
rect 1500 -1720 1700 -1520
rect 3584 -1946 3784 -1940
rect 3584 -2134 3590 -1946
rect 3590 -2134 3778 -1946
rect 3778 -2134 3784 -1946
rect 3584 -2140 3784 -2134
rect 3194 -2460 3394 -2260
rect 1500 -3080 1700 -2880
rect 1110 -3590 1310 -3390
rect 1500 -3396 1700 -3390
rect 1500 -3584 1506 -3396
rect 1506 -3584 1694 -3396
rect 1694 -3584 1700 -3396
rect 1500 -3590 1700 -3584
rect 2240 -3587 2294 -3443
rect 2432 -3587 2486 -3443
rect 2624 -3587 2678 -3443
rect 2816 -3587 2870 -3443
rect 3008 -3587 3062 -3443
rect 2336 -4219 2390 -4075
rect 2528 -4219 2582 -4075
rect 2720 -4219 2774 -4075
rect 2912 -4219 2966 -4075
rect 4704 -2460 4904 -2260
rect 3964 -3026 4164 -3020
rect 3964 -3214 3970 -3026
rect 3970 -3214 4158 -3026
rect 4158 -3214 4164 -3026
rect 3964 -3220 4164 -3214
rect 3584 -3590 3784 -3390
rect 1500 -4690 1700 -4490
rect 3196 -4890 3396 -4690
rect 2242 -5076 2296 -4932
rect 2434 -5076 2488 -4932
rect 2626 -5076 2680 -4932
rect 2818 -5076 2872 -4932
rect 3010 -5076 3064 -4932
rect 2338 -5708 2392 -5564
rect 2530 -5708 2584 -5564
rect 2722 -5708 2776 -5564
rect 2914 -5708 2968 -5564
rect 5358 -3660 5558 -3460
rect 4504 -4570 4704 -4370
rect 3994 -5076 4048 -4932
rect 4186 -5076 4240 -4932
rect 4378 -5076 4432 -4932
rect 4570 -5076 4624 -4932
rect 4762 -5076 4816 -4932
rect 4090 -5708 4144 -5564
rect 4282 -5708 4336 -5564
rect 4474 -5708 4528 -5564
rect 4666 -5708 4720 -5564
rect 5358 -5566 5558 -5560
rect 5358 -5754 5364 -5566
rect 5364 -5754 5552 -5566
rect 5552 -5754 5558 -5566
rect 5358 -5760 5558 -5754
rect 1500 -6180 1700 -5980
<< metal2 >>
rect 1500 -1520 1700 -1514
rect 1700 -1720 2650 -1520
rect 1500 -1726 1700 -1720
rect 1910 -2140 2110 -1940
rect 710 -2460 2110 -2260
rect 2450 -2460 2650 -1720
rect 3584 -1940 3784 -1934
rect 3784 -2140 4154 -1940
rect 3584 -2146 3784 -2140
rect 3194 -2260 3394 -2254
rect 3394 -2460 4164 -2260
rect 4504 -2460 4704 -2260
rect 4904 -2460 4910 -2260
rect 3194 -2466 3394 -2460
rect 1500 -2880 1700 -2874
rect 710 -3080 1500 -2880
rect 1500 -3086 1700 -3080
rect 1910 -3020 2110 -2570
rect 3194 -2770 4164 -2570
rect 3194 -3020 3394 -2770
rect 1910 -3220 3394 -3020
rect 3964 -3020 4164 -2770
rect 1110 -3390 1310 -3384
rect 710 -3590 1110 -3390
rect 1310 -3590 1500 -3390
rect 1700 -3443 3584 -3390
rect 1700 -3587 2240 -3443
rect 2294 -3587 2432 -3443
rect 2486 -3587 2624 -3443
rect 2678 -3587 2816 -3443
rect 2870 -3587 3008 -3443
rect 3062 -3587 3584 -3443
rect 1700 -3590 3584 -3587
rect 3784 -3590 3790 -3390
rect 3964 -3460 4164 -3220
rect 5358 -3460 5558 -3454
rect 1110 -3596 1310 -3590
rect 3964 -3660 5358 -3460
rect 5358 -3666 5558 -3660
rect 1500 -4075 3080 -4070
rect 1500 -4130 2336 -4075
rect 710 -4219 2336 -4130
rect 2390 -4219 2528 -4075
rect 2582 -4219 2720 -4075
rect 2774 -4219 2912 -4075
rect 2966 -4219 3080 -4075
rect 710 -4270 3080 -4219
rect 710 -4330 1700 -4270
rect 710 -4690 1500 -4490
rect 1700 -4690 1706 -4490
rect 3196 -4570 4504 -4370
rect 4704 -4570 4710 -4370
rect 3196 -4690 3396 -4570
rect 1810 -4932 3080 -4880
rect 3190 -4890 3196 -4690
rect 3396 -4890 3402 -4690
rect 1810 -5076 2242 -4932
rect 2296 -5076 2434 -4932
rect 2488 -5076 2626 -4932
rect 2680 -5076 2818 -4932
rect 2872 -5076 3010 -4932
rect 3064 -5076 3080 -4932
rect 1810 -5080 3080 -5076
rect 3984 -4932 5958 -4880
rect 3984 -5076 3994 -4932
rect 4048 -5076 4186 -4932
rect 4240 -5076 4378 -4932
rect 4432 -5076 4570 -4932
rect 4624 -5076 4762 -4932
rect 4816 -5076 5958 -4932
rect 3984 -5080 5958 -5076
rect 1810 -5280 2010 -5080
rect 710 -5480 2010 -5280
rect 1500 -5564 5358 -5560
rect 1500 -5620 2338 -5564
rect 710 -5708 2338 -5620
rect 2392 -5708 2530 -5564
rect 2584 -5708 2722 -5564
rect 2776 -5708 2914 -5564
rect 2968 -5708 4090 -5564
rect 4144 -5708 4282 -5564
rect 4336 -5708 4474 -5564
rect 4528 -5708 4666 -5564
rect 4720 -5708 5358 -5564
rect 710 -5760 5358 -5708
rect 5558 -5760 5564 -5560
rect 710 -5820 1700 -5760
rect 710 -6180 1500 -5980
rect 1700 -6180 1706 -5980
use level_shifter_dd  level_shifter_dd_0
timestamp 1713791489
transform 1 0 1690 0 1 -1070
box 220 -1910 960 -652
use level_shifter_dd  level_shifter_dd_1
timestamp 1713791489
transform 1 0 3744 0 1 -1070
box 220 -1910 960 -652
use sky130_fd_pr__nfet_01v8_HNLS5R  sky130_fd_pr__nfet_01v8_HNLS5R_0
timestamp 1713791489
transform 1 0 4405 0 1 -5320
box -551 -610 551 610
use sky130_fd_pr__pfet_01v8_XGNZDL  sky130_fd_pr__pfet_01v8_XGNZDL_0
timestamp 1713791715
transform 1 0 2651 0 1 -3831
box -551 -619 551 619
use sky130_fd_pr__nfet_01v8_HNLS5R  XM18
timestamp 1713791489
transform 1 0 2653 0 1 -5320
box -551 -610 551 610
<< labels >>
flabel metal2 710 -2460 910 -2260 0 FreeSans 256 0 0 0 ENA
port 2 nsew
flabel metal2 710 -3080 910 -2880 0 FreeSans 256 0 0 0 ENA_B
port 3 nsew
flabel metal2 710 -3590 910 -3390 0 FreeSans 256 0 0 0 DVDD
port 1 nsew
flabel metal2 710 -4690 910 -4490 0 FreeSans 256 0 0 0 STDBY
port 4 nsew
flabel metal2 710 -4330 910 -4130 0 FreeSans 256 0 0 0 SG_DVDD
port 7 nsew
flabel metal2 710 -6180 910 -5980 0 FreeSans 256 0 0 0 STDBY_B
port 5 nsew
flabel metal2 710 -5480 910 -5280 0 FreeSans 256 0 0 0 SG_DVSS
port 6 nsew
flabel metal2 710 -5820 910 -5620 0 FreeSans 256 0 0 0 DVSS
port 0 nsew
flabel metal2 5758 -5080 5958 -4880 0 FreeSans 256 0 0 0 DOUT
port 8 nsew
<< end >>
