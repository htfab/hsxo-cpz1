magic
tech sky130A
magscale 1 2
timestamp 1713795963
<< error_s >>
rect 3828 11829 3862 12212
rect 3950 11889 4008 11903
rect 4108 11889 4166 11903
rect 4024 11849 4092 11863
rect 3896 11835 4220 11849
rect 4008 11829 4130 11835
rect 4254 11829 4288 12212
rect 4438 11829 4472 12212
rect 4560 11889 4618 11903
rect 4718 11889 4776 11903
rect 4634 11849 4702 11863
rect 4506 11835 4830 11849
rect 4618 11829 4740 11835
rect 4864 11829 4898 12212
rect 4967 11829 5432 11938
rect 6711 11829 7174 11938
rect 7248 11829 7282 12212
rect 7370 11889 7428 11903
rect 7528 11889 7586 11903
rect 7444 11849 7512 11863
rect 7316 11835 7640 11849
rect 7428 11829 7550 11835
rect 7674 11829 7708 12212
rect 7858 11829 7892 12212
rect 7980 11889 8038 11903
rect 8138 11889 8196 11903
rect 8054 11849 8122 11863
rect 7926 11835 8250 11849
rect 8038 11829 8160 11835
rect 8284 11829 8318 12212
rect 2667 11795 8693 11829
rect 3828 11766 3862 11795
rect 4008 11792 4108 11795
rect 4254 11766 4288 11795
rect 4438 11766 4472 11795
rect 4618 11792 4718 11795
rect 4864 11766 4898 11795
rect 4967 11730 5432 11795
rect 4852 11716 5432 11730
rect 4967 11702 5432 11716
rect 4880 11688 5432 11702
rect 4967 11542 5432 11688
rect 6711 11736 7174 11795
rect 7248 11766 7282 11795
rect 7428 11792 7528 11795
rect 7674 11766 7708 11795
rect 7858 11766 7892 11795
rect 8038 11792 8138 11795
rect 8284 11766 8318 11795
rect 6711 11730 7218 11736
rect 6711 11716 7298 11730
rect 6711 11708 7174 11716
rect 6711 11702 7190 11708
rect 6711 11688 7270 11702
rect 6711 11542 7174 11688
rect 8719 11542 8753 11769
rect 3990 11538 4730 11542
rect 3780 11186 4946 11538
rect 4950 11186 7190 11542
rect 7410 11538 8160 11542
rect 8360 11538 8840 11542
rect 7111 11142 7174 11186
rect 7184 10906 7190 11186
rect 7111 10822 7190 10906
rect 7200 10822 8840 11538
rect 7171 10768 7184 10822
rect 7170 10368 7184 10560
rect 8719 7828 8753 10822
rect 7744 7794 9118 7828
rect 8719 7728 8753 7794
rect 8702 7717 8753 7728
rect 8699 7690 8753 7717
rect 8754 7690 8773 7728
rect 8685 7663 8753 7690
rect 8765 7663 8773 7690
rect 8685 7656 8773 7663
rect 8776 7656 8787 7690
rect 8792 7656 8811 7690
rect 8699 7631 8718 7656
rect 8719 7631 8773 7656
rect 8696 7597 8773 7631
rect 8699 6821 8787 7597
rect 8984 7012 9040 7016
rect 8840 6972 9046 7012
rect 8840 6956 9096 6972
rect 8699 6809 8773 6821
rect 8840 6812 9040 6956
rect 8699 6800 8718 6809
rect 8719 6800 8753 6809
rect 8765 6800 8773 6809
rect 8699 6762 8753 6800
rect 8754 6762 8773 6800
rect 8685 6728 8753 6762
rect 8699 6712 8718 6728
rect 8699 6701 8710 6712
rect 8719 6624 8753 6728
rect 8765 6701 8773 6762
rect 8776 6728 8787 6762
rect 8792 6728 8811 6762
rect 7744 6590 9118 6624
rect 8719 6502 8753 6590
rect 8670 4906 8840 6502
rect 9224 6472 9280 6528
rect 9280 6416 9336 6472
rect 8830 3336 8838 3338
rect 8802 3308 8810 3310
rect 3900 3012 4646 3156
rect 3735 2971 4646 3012
rect 3735 2954 5188 2971
rect 3900 2942 5188 2954
rect 5290 2942 7600 3156
rect 3900 2868 7600 2942
rect 3760 2648 7600 2868
rect 3937 2602 4011 2648
rect 4026 2604 7600 2648
rect 4026 2602 4246 2604
rect 3760 2382 4246 2602
rect 4360 2477 7306 2604
rect 3900 2296 4186 2382
rect 4332 2312 7306 2477
rect 4332 2296 5173 2312
rect 3735 2279 5173 2296
rect 3735 2238 4646 2279
rect 3900 1982 4186 2238
rect 4360 1982 4646 2238
rect 4916 2078 4920 2279
rect 4944 2112 4948 2242
rect 4950 2241 5150 2279
rect 4950 2112 5156 2241
rect 5000 2082 5080 2112
rect 5132 2106 5150 2112
rect 5160 2084 5184 2241
rect 5311 2123 7306 2312
rect 5160 2078 5178 2084
rect 1740 1456 1940 1458
rect 1740 1312 1940 1452
rect 1740 1252 2100 1312
rect 1900 1112 2100 1252
rect 4360 -118 4440 1982
rect 7174 1972 7306 2123
rect 7314 2123 7600 2604
rect 8802 3144 8814 3308
rect 8802 2510 8810 3144
rect 8830 3116 8842 3336
rect 9274 3168 9330 3196
rect 9243 3142 9330 3168
rect 8830 2482 8838 3116
rect 9271 3114 9330 3140
rect 9274 3086 9330 3114
rect 7676 2346 7734 2427
rect 7676 2288 7765 2346
rect 7314 1972 7560 2123
rect 7314 1832 7446 1972
rect 9980 1682 10780 2482
rect 8802 -120 8920 -111
rect 7492 -138 8920 -120
rect 8830 -148 8948 -139
rect 7520 -166 8948 -148
rect 7314 -760 7520 -288
rect 7314 -818 7534 -760
rect 4662 -1013 7534 -818
rect 4662 -1104 7520 -1013
rect 7892 -1400 8320 -1394
rect 3842 -1404 8320 -1400
rect 7920 -1428 8320 -1422
rect 3870 -1432 8320 -1428
<< metal1 >>
rect 0 16110 30870 16310
rect 31070 16110 31076 16310
rect 0 602 200 16110
rect 8834 14970 8840 15170
rect 9040 14970 24190 15170
rect 24390 14970 24396 15170
rect 9704 9950 9710 10150
rect 9910 9950 9916 10150
rect 744 9510 750 9710
rect 950 9510 956 9710
rect 364 7042 370 7250
rect 570 7042 576 7250
rect -6 400 0 602
rect 200 400 206 602
rect 370 -6750 570 7042
rect 750 5572 950 9510
rect 8840 7012 9040 7018
rect 9710 7012 9910 9950
rect 9040 6812 9910 7012
rect 8840 6806 9040 6812
rect 8834 6390 8840 6590
rect 9040 6390 9480 6590
rect 8824 6000 8830 6200
rect 9030 6000 9036 6200
rect 744 5372 750 5572
rect 950 5372 956 5572
rect 1124 -348 1130 -148
rect 1330 -348 1336 -148
rect 1130 -6340 1330 -348
rect 8830 -630 9030 6000
rect 8824 -830 8830 -630
rect 9030 -830 9036 -630
rect 9280 -680 9480 6390
rect 9280 -880 9710 -680
rect 9910 -880 9916 -680
rect 30870 -4510 31070 -4504
rect 30870 -6340 31070 -4710
rect 1130 -6540 31070 -6340
rect 370 -6950 19620 -6750
rect 19820 -6950 19826 -6750
<< via1 >>
rect 30870 16110 31070 16310
rect 8840 14970 9040 15170
rect 24190 14970 24390 15170
rect 9710 9950 9910 10150
rect 750 9510 950 9710
rect 370 7042 570 7250
rect 0 400 200 602
rect 8840 6812 9040 7012
rect 8840 6390 9040 6590
rect 8830 6000 9030 6200
rect 750 5372 950 5572
rect 1130 -348 1330 -148
rect 8830 -830 9030 -630
rect 9710 -880 9910 -680
rect 30870 -4710 31070 -4510
rect 19620 -6950 19820 -6750
<< metal2 >>
rect 30870 16310 31070 16316
rect 0 16305 200 16310
rect -4 16115 5 16305
rect 195 16115 204 16305
rect 0 6860 200 16115
rect 370 16110 9480 16310
rect 370 9280 570 16110
rect 8840 15170 9040 15176
rect 1121 11302 1130 11502
rect 1330 11302 1339 11502
rect 750 9710 950 9716
rect 741 9510 750 9710
rect 950 9510 959 9710
rect 750 9504 950 9510
rect 370 9080 950 9280
rect 370 7250 570 7256
rect 361 7050 370 7250
rect 570 7050 579 7250
rect 366 7047 370 7050
rect 570 7047 574 7050
rect 370 7036 570 7042
rect 0 6651 200 6660
rect 750 5977 950 9080
rect 1121 7442 1130 7642
rect 1330 7442 1339 7642
rect 1121 7042 1130 7242
rect 1330 7042 1339 7242
rect 8840 7172 9040 14970
rect 8834 6812 8840 7012
rect 9040 6812 9046 7012
rect 8840 6590 9040 6596
rect 8840 6384 9040 6390
rect 8830 6200 9030 6206
rect 8830 5994 9030 6000
rect 750 5787 755 5977
rect 945 5787 950 5977
rect 750 5782 950 5787
rect 1121 5782 1130 5982
rect 1330 5782 1339 5982
rect 755 5778 945 5782
rect 750 5572 950 5578
rect 950 5372 1330 5572
rect 9280 5380 9480 16110
rect 25870 16050 26070 16059
rect 30870 15900 31070 16110
rect 24190 15170 24390 15176
rect 9710 10150 9910 10156
rect 24190 9950 24390 14970
rect 9710 9944 9910 9950
rect 25870 6270 26070 15850
rect 24200 6070 26070 6270
rect 750 5366 950 5372
rect 9280 5180 9910 5380
rect 9271 2940 9280 3140
rect 9480 2940 9910 3140
rect 1121 1872 1130 2072
rect 1330 1872 1339 2072
rect 730 1550 930 1559
rect 0 602 200 608
rect -9 400 0 600
rect 200 400 209 600
rect 0 394 200 400
rect 730 237 930 1350
rect 1121 742 1130 942
rect 1330 742 1339 942
rect 1121 402 1130 602
rect 1330 402 1339 602
rect 730 47 735 237
rect 925 47 930 237
rect 730 42 930 47
rect 1121 42 1130 242
rect 1330 42 1339 242
rect 27640 100 27980 300
rect 735 38 925 42
rect 1130 -148 1330 -142
rect 1130 -354 1330 -348
rect 8830 -148 9030 -139
rect 8830 -357 9030 -348
rect 1121 -688 1130 -488
rect 1330 -688 1339 -488
rect 8830 -630 9030 -624
rect 8830 -6340 9030 -830
rect 9710 -680 9910 -674
rect 9710 -886 9910 -880
rect 19155 -6340 19345 -6336
rect 8830 -6345 19350 -6340
rect 8830 -6535 19155 -6345
rect 19345 -6535 19350 -6345
rect 8830 -6540 19350 -6535
rect 19155 -6544 19345 -6540
rect 19620 -6750 19820 -5920
rect 24210 -6340 24410 -4320
rect 27640 -4510 27840 100
rect 30864 -4710 30870 -4510
rect 31070 -4710 31076 -4510
rect 27640 -4719 27840 -4710
rect 20091 -6540 20100 -6340
rect 20300 -6540 24410 -6340
rect 31540 -6750 31740 300
rect 31531 -6950 31540 -6750
rect 31740 -6950 31749 -6750
rect 19620 -6956 19820 -6950
<< via2 >>
rect 5 16115 195 16305
rect 1130 11302 1330 11502
rect 750 9510 950 9710
rect 370 7050 570 7250
rect 375 7047 565 7050
rect 0 6660 200 6860
rect 1130 7442 1330 7642
rect 1130 7042 1330 7242
rect 755 5787 945 5977
rect 1130 5782 1330 5982
rect 25870 15850 26070 16050
rect 9280 2940 9480 3140
rect 1130 1872 1330 2072
rect 730 1350 930 1550
rect 0 400 200 600
rect 1130 742 1330 942
rect 1130 402 1330 602
rect 735 47 925 237
rect 1130 42 1330 242
rect 8830 -348 9030 -148
rect 1130 -688 1330 -488
rect 19155 -6535 19345 -6345
rect 27640 -4710 27840 -4510
rect 20100 -6540 20300 -6340
rect 31540 -6950 31740 -6750
<< metal3 >>
rect 0 16305 9480 16310
rect 0 16115 5 16305
rect 195 16115 9480 16305
rect 0 16110 9480 16115
rect 1125 11502 1335 11507
rect -200 11302 1130 11502
rect 1330 11302 1335 11502
rect -200 11300 0 11302
rect 1125 11297 1335 11302
rect 745 9710 955 9715
rect -200 9510 750 9710
rect 950 9510 955 9710
rect 745 9505 955 9510
rect 1125 7642 1335 7647
rect -200 7442 1130 7642
rect 1330 7442 1335 7642
rect -200 7440 0 7442
rect 1125 7437 1335 7442
rect 365 7250 575 7255
rect 365 7050 370 7250
rect 570 7242 575 7250
rect 1125 7242 1335 7247
rect 570 7050 1130 7242
rect 365 7047 375 7050
rect 565 7047 1130 7050
rect 365 7045 1130 7047
rect 370 7042 1130 7045
rect 1330 7042 1335 7242
rect 1125 7037 1335 7042
rect -5 6860 205 6865
rect -200 6660 0 6860
rect 200 6660 205 6860
rect -5 6655 205 6660
rect 1125 5982 1335 5987
rect -200 5977 1130 5982
rect -200 5787 755 5977
rect 945 5787 1130 5977
rect -200 5782 1130 5787
rect 1330 5782 1335 5982
rect -200 5780 0 5782
rect 1125 5777 1335 5782
rect 9280 3145 9480 16110
rect 25865 16050 26075 16055
rect 25865 16045 25870 16050
rect 26070 16045 26075 16050
rect 25865 15839 26075 15845
rect 9275 3140 9485 3145
rect 9275 2940 9280 3140
rect 9480 2940 9485 3140
rect 9275 2935 9485 2940
rect 1125 2072 1335 2077
rect -200 1872 1130 2072
rect 1330 1872 1335 2072
rect -200 1870 0 1872
rect 1125 1867 1335 1872
rect 725 1550 935 1555
rect -200 1350 730 1550
rect 930 1350 935 1550
rect 725 1345 935 1350
rect 1125 942 1335 947
rect -200 742 1130 942
rect 1330 742 1335 942
rect -200 740 0 742
rect 1125 737 1335 742
rect -5 602 205 605
rect 1125 602 1335 607
rect -5 600 1130 602
rect -5 400 0 600
rect 200 402 1130 600
rect 1330 402 1335 602
rect 200 400 205 402
rect -5 395 205 400
rect 1125 397 1335 402
rect 1125 242 1335 247
rect 730 237 1130 242
rect 730 47 735 237
rect 925 47 1130 237
rect 730 42 1130 47
rect 1330 42 1335 242
rect 1125 37 1335 42
rect 8825 -148 9035 -143
rect 8825 -348 8830 -148
rect 9030 -348 9035 -148
rect 8825 -353 9035 -348
rect 1125 -488 1335 -483
rect -200 -688 1130 -488
rect 1330 -688 1335 -488
rect -200 -690 0 -688
rect 1125 -693 1335 -688
rect 8830 -6750 9030 -353
rect 27635 -4505 27845 -4499
rect 27635 -4710 27640 -4705
rect 27840 -4710 27845 -4705
rect 27635 -4715 27845 -4710
rect 20095 -6340 20305 -6335
rect 19150 -6345 20100 -6340
rect 19150 -6535 19155 -6345
rect 19345 -6535 20100 -6345
rect 19150 -6540 20100 -6535
rect 20300 -6540 20305 -6340
rect 20095 -6545 20305 -6540
rect 31535 -6750 31745 -6745
rect 8830 -6950 31540 -6750
rect 31740 -6950 31950 -6750
rect 31535 -6955 31745 -6950
<< via3 >>
rect 25865 15850 25870 16045
rect 25870 15850 26070 16045
rect 26070 15850 26075 16045
rect 25865 15845 26075 15850
rect 27635 -4510 27845 -4505
rect 27635 -4705 27640 -4510
rect 27640 -4705 27840 -4510
rect 27840 -4705 27845 -4510
<< metal4 >>
rect 25864 16045 26076 16046
rect 25864 15845 25865 16045
rect 26075 15845 26076 16045
rect 25864 15844 26076 15845
rect 25870 -4260 26070 15844
rect 27640 -4504 27840 15660
rect 27634 -4505 27846 -4504
rect 27634 -4705 27635 -4505
rect 27845 -4705 27846 -4505
rect 27634 -4706 27846 -4705
use power_gating  power_gating_0
timestamp 1713795963
transform 1 0 1870 0 1 10256
box -834 -14876 9710 5689
use schmitt_trigger_pullmid  schmitt_trigger_pullmid_0
timestamp 1713748097
transform 1 0 26390 0 1 -720
box 1390 -3990 5350 16820
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  sky130_fd_pr__cap_mim_m3_1_MPZGNS_0
timestamp 1713748097
transform 1 0 26106 0 1 5700
box -1686 -9960 1686 9960
use vittoz_pierce_osc  vittoz_pierce_osc_0
timestamp 1713748602
transform 1 0 10050 0 1 -2190
box -340 -3940 14370 18841
<< labels >>
flabel metal3 -200 11300 0 11500 0 FreeSans 256 0 0 0 AVDD
port 5 nsew
flabel metal3 -200 9510 0 9710 0 FreeSans 256 0 0 0 AVSS
port 7 nsew
flabel metal3 -200 7440 0 7640 0 FreeSans 256 0 0 0 IBIAS
port 9 nsew
flabel metal3 -200 6660 0 6860 0 FreeSans 256 0 0 0 XOUT
port 0 nsew
flabel metal3 -200 5780 0 5980 0 FreeSans 256 0 0 0 XIN
port 1 nsew
flabel metal3 -200 1870 0 2070 0 FreeSans 256 0 0 0 ENA
port 2 nsew
flabel metal3 -200 1350 0 1550 0 FreeSans 256 0 0 0 STDBY
port 3 nsew
flabel metal3 -200 740 0 940 0 FreeSans 256 0 0 0 DVDD
port 6 nsew
flabel metal3 -200 -690 0 -490 0 FreeSans 256 0 0 0 DVSS
port 8 nsew
flabel metal3 31750 -6950 31950 -6750 0 FreeSans 256 0 0 0 DOUT
port 4 nsew
<< end >>
