magic
tech sky130A
magscale 1 2
timestamp 1718125978
<< pwell >>
rect -782 -2182 782 2182
<< psubdiff >>
rect -746 2112 -650 2146
rect 650 2112 746 2146
rect -746 2050 -712 2112
rect 712 2050 746 2112
rect -746 -2112 -712 -2050
rect 712 -2112 746 -2050
rect -746 -2146 -650 -2112
rect 650 -2146 746 -2112
<< psubdiffcont >>
rect -650 2112 650 2146
rect -746 -2050 -712 2050
rect 712 -2050 746 2050
rect -650 -2146 650 -2112
<< xpolycontact >>
rect -616 1584 -546 2016
rect -616 -2016 -546 -1584
rect -450 1584 -380 2016
rect -450 -2016 -380 -1584
rect -284 1584 -214 2016
rect -284 -2016 -214 -1584
rect -118 1584 -48 2016
rect -118 -2016 -48 -1584
rect 48 1584 118 2016
rect 48 -2016 118 -1584
rect 214 1584 284 2016
rect 214 -2016 284 -1584
rect 380 1584 450 2016
rect 380 -2016 450 -1584
rect 546 1584 616 2016
rect 546 -2016 616 -1584
<< xpolyres >>
rect -616 -1584 -546 1584
rect -450 -1584 -380 1584
rect -284 -1584 -214 1584
rect -118 -1584 -48 1584
rect 48 -1584 118 1584
rect 214 -1584 284 1584
rect 380 -1584 450 1584
rect 546 -1584 616 1584
<< locali >>
rect -746 2112 -650 2146
rect 650 2112 746 2146
rect -746 2050 -712 2112
rect 712 2050 746 2112
rect -746 -2112 -712 -2050
rect 712 -2112 746 -2050
rect -746 -2146 -650 -2112
rect 650 -2146 746 -2112
<< viali >>
rect -600 1601 -562 1998
rect -434 1601 -396 1998
rect -268 1601 -230 1998
rect -102 1601 -64 1998
rect 64 1601 102 1998
rect 230 1601 268 1998
rect 396 1601 434 1998
rect 562 1601 600 1998
rect -600 -1998 -562 -1601
rect -434 -1998 -396 -1601
rect -268 -1998 -230 -1601
rect -102 -1998 -64 -1601
rect 64 -1998 102 -1601
rect 230 -1998 268 -1601
rect 396 -1998 434 -1601
rect 562 -1998 600 -1601
<< metal1 >>
rect -606 1998 -556 2010
rect -606 1601 -600 1998
rect -562 1601 -556 1998
rect -606 1589 -556 1601
rect -440 1998 -390 2010
rect -440 1601 -434 1998
rect -396 1601 -390 1998
rect -440 1589 -390 1601
rect -274 1998 -224 2010
rect -274 1601 -268 1998
rect -230 1601 -224 1998
rect -274 1589 -224 1601
rect -108 1998 -58 2010
rect -108 1601 -102 1998
rect -64 1601 -58 1998
rect -108 1589 -58 1601
rect 58 1998 108 2010
rect 58 1601 64 1998
rect 102 1601 108 1998
rect 58 1589 108 1601
rect 224 1998 274 2010
rect 224 1601 230 1998
rect 268 1601 274 1998
rect 224 1589 274 1601
rect 390 1998 440 2010
rect 390 1601 396 1998
rect 434 1601 440 1998
rect 390 1589 440 1601
rect 556 1998 606 2010
rect 556 1601 562 1998
rect 600 1601 606 1998
rect 556 1589 606 1601
rect -606 -1601 -556 -1589
rect -606 -1998 -600 -1601
rect -562 -1998 -556 -1601
rect -606 -2010 -556 -1998
rect -440 -1601 -390 -1589
rect -440 -1998 -434 -1601
rect -396 -1998 -390 -1601
rect -440 -2010 -390 -1998
rect -274 -1601 -224 -1589
rect -274 -1998 -268 -1601
rect -230 -1998 -224 -1601
rect -274 -2010 -224 -1998
rect -108 -1601 -58 -1589
rect -108 -1998 -102 -1601
rect -64 -1998 -58 -1601
rect -108 -2010 -58 -1998
rect 58 -1601 108 -1589
rect 58 -1998 64 -1601
rect 102 -1998 108 -1601
rect 58 -2010 108 -1998
rect 224 -1601 274 -1589
rect 224 -1998 230 -1601
rect 268 -1998 274 -1601
rect 224 -2010 274 -1998
rect 390 -1601 440 -1589
rect 390 -1998 396 -1601
rect 434 -1998 440 -1601
rect 390 -2010 440 -1998
rect 556 -1601 606 -1589
rect 556 -1998 562 -1601
rect 600 -1998 606 -1601
rect 556 -2010 606 -1998
<< properties >>
string FIXED_BBOX -729 -2129 729 2129
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 16 m 1 nx 8 wmin 0.350 lmin 0.50 rho 2000 val 92.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
