magic
tech sky130A
magscale 1 2
timestamp 1713816941
<< mvpsubdiff >>
rect -87 15225 -63 15259
rect 7043 15225 7067 15259
rect -523 14799 -489 14823
rect -523 3059 -489 3083
rect 7469 14799 7503 14823
rect 10443 13449 10467 13483
rect 19883 13449 19907 13483
rect 21193 13449 21217 13483
rect 23453 13449 23477 13483
rect 7469 3059 7503 3083
rect 10007 13023 10041 13047
rect -87 2623 -63 2657
rect 7043 2623 7067 2657
rect -637 1335 -613 1369
rect 4053 1335 4077 1369
rect -1073 909 -1039 933
rect -1073 -4341 -1039 -4317
rect 4479 909 4513 933
rect 10007 -1847 10041 -1823
rect 20309 13023 20343 13047
rect 20757 13023 20791 13047
rect 20757 2583 20791 2607
rect 23879 13023 23913 13047
rect 28074 3708 28098 3742
rect 31432 3708 31456 3742
rect 23879 2583 23913 2607
rect 27638 3282 27672 3306
rect 21193 2147 21217 2181
rect 23453 2147 23477 2181
rect 20309 -1847 20343 -1823
rect 10443 -2283 10467 -2249
rect 19883 -2283 19907 -2249
rect 27638 -2876 27672 -2852
rect 31858 3282 31892 3306
rect 31858 -2876 31892 -2852
rect 28074 -3312 28098 -3278
rect 31432 -3312 31456 -3278
rect 4479 -4341 4513 -4317
rect -637 -4777 -613 -4743
rect 4053 -4777 4077 -4743
<< mvpsubdiffcont >>
rect -63 15225 7043 15259
rect -523 3083 -489 14799
rect 7469 3083 7503 14799
rect 10467 13449 19883 13483
rect 21217 13449 23453 13483
rect -63 2623 7043 2657
rect -613 1335 4053 1369
rect -1073 -4317 -1039 909
rect 4479 -4317 4513 909
rect 10007 -1823 10041 13023
rect 20309 -1823 20343 13023
rect 20757 2607 20791 13023
rect 23879 2607 23913 13023
rect 28098 3708 31432 3742
rect 21217 2147 23453 2181
rect 10467 -2283 19883 -2249
rect 27638 -2852 27672 3282
rect 31858 -2852 31892 3282
rect 28098 -3312 31432 -3278
rect -613 -4777 4053 -4743
<< locali >>
rect -1670 15259 32490 15870
rect -1670 15225 -63 15259
rect 7043 15225 32490 15259
rect -1670 15070 32490 15225
rect -1673 15025 32490 15070
rect -1673 14799 -289 15025
rect -1673 3083 -523 14799
rect -489 3083 -289 14799
rect -1673 2857 -289 3083
rect 7269 14799 32490 15025
rect 7269 3083 7469 14799
rect 7503 13483 32490 14799
rect 7503 13449 10467 13483
rect 19883 13449 21217 13483
rect 23453 13449 32490 13483
rect 7503 13249 32490 13449
rect 7503 13023 10241 13249
rect 7503 3083 10007 13023
rect 7269 2857 10007 3083
rect -1673 2657 10007 2857
rect -1673 2623 -63 2657
rect 7043 2623 10007 2657
rect -1673 1369 10007 2623
rect -1673 1335 -613 1369
rect 4053 1335 10007 1369
rect -1673 1135 10007 1335
rect -1673 909 -839 1135
rect -1673 -4317 -1073 909
rect -1039 -4317 -839 909
rect -1673 -4543 -839 -4317
rect 4279 909 10007 1135
rect 4279 -4317 4479 909
rect 4513 -1823 10007 909
rect 10041 -1823 10241 13023
rect 4513 -2049 10241 -1823
rect 20109 13023 20991 13249
rect 20109 -1823 20309 13023
rect 20343 2607 20757 13023
rect 20791 2607 20991 13023
rect 20343 2381 20991 2607
rect 23679 13023 32490 13249
rect 23679 2607 23879 13023
rect 23913 4342 32490 13023
rect 23913 3742 32492 4342
rect 23913 3708 28098 3742
rect 31432 3708 32492 3742
rect 23913 3508 32492 3708
rect 23913 3282 27872 3508
rect 23913 2607 27638 3282
rect 23679 2381 27638 2607
rect 20343 2181 27638 2381
rect 20343 2147 21217 2181
rect 23453 2147 27638 2181
rect 20343 -1823 27638 2147
rect 20109 -2049 27638 -1823
rect 4513 -2249 27638 -2049
rect 4513 -2283 10467 -2249
rect 19883 -2283 27638 -2249
rect 4513 -2852 27638 -2283
rect 27672 -2852 27872 3282
rect 4513 -3078 27872 -2852
rect 31658 3282 32492 3508
rect 31658 -2852 31858 3282
rect 31892 -2852 32490 3282
rect 31658 -3078 32492 -2852
rect 4513 -3278 32492 -3078
rect 4513 -3312 28098 -3278
rect 31432 -3312 32492 -3278
rect 4513 -3912 32492 -3312
rect 4513 -4317 32490 -3912
rect 4279 -4543 32490 -4317
rect -1673 -4577 32490 -4543
rect -2346 -4743 32490 -4577
rect -2346 -4777 -613 -4743
rect 4053 -4777 32490 -4743
rect -2346 -5377 32490 -4777
rect 4700 -5380 32490 -5377
<< viali >>
rect -3146 -5377 -2346 -4577
<< metal1 >>
rect 2114 17740 2914 17746
rect 2108 17734 2920 17740
rect 2108 16940 2114 17734
rect 2914 16940 2920 17734
rect 7964 17090 7970 17490
rect 8370 17090 8376 17490
rect 2114 16928 2914 16934
rect 2414 14888 2614 16928
rect -396 2300 -196 2700
rect 24 2696 224 2702
rect 24 2490 224 2496
rect -396 2100 5620 2300
rect 4784 -2814 4790 -2414
rect 5190 -2814 5196 -2414
rect 5420 -2690 5620 2100
rect 7970 -1824 8370 17090
rect 22820 16720 23620 16726
rect 8760 15920 22820 16720
rect 23620 15920 23630 16720
rect 8760 12340 9560 15920
rect 22820 15914 23620 15920
rect 8760 11534 9560 11540
rect 8754 9950 8760 10750
rect 9560 9950 9566 10750
rect 8760 7492 9560 9950
rect 8754 6692 8760 7492
rect 9560 6692 9566 7492
rect 8754 5416 8760 6216
rect 9560 5416 9566 6216
rect 8760 -80 9560 5416
rect 8754 -880 8760 -80
rect 9560 -880 9566 -80
rect 7964 -2224 7970 -1824
rect 8370 -2224 8376 -1824
rect 4364 -3234 4370 -3034
rect 4570 -3234 4576 -3034
rect 4790 -3170 5190 -2814
rect 5420 -2890 9020 -2690
rect 4370 -3880 4570 -3234
rect 4790 -3570 7960 -3170
rect 4370 -4080 7280 -3880
rect -3152 -4571 -2340 -4565
rect -3158 -5383 -3152 -4571
rect -2352 -4577 -2340 -4571
rect -2346 -5377 -2340 -4577
rect -2352 -5383 -2340 -5377
rect -3152 -5389 -2340 -5383
rect 7080 -6770 7280 -4080
rect 7560 -6090 7960 -3570
rect 8820 -5530 9020 -2890
rect 19620 -5530 19820 -5220
rect 8820 -5730 19820 -5530
rect 7560 -6490 30770 -6090
rect 31170 -6490 31176 -6090
rect 31545 -6510 32345 -6504
rect 31530 -6770 31545 -6510
rect 7080 -6970 31545 -6770
rect 31530 -7110 31545 -6970
rect 31530 -7310 31540 -7110
rect 31540 -7316 32345 -7310
<< via1 >>
rect 2114 16934 2914 17734
rect 7970 17090 8370 17490
rect 24 2496 224 2696
rect 4790 -2814 5190 -2414
rect 22820 15920 23620 16720
rect 8760 11540 9560 12340
rect 8760 9950 9560 10750
rect 8760 6692 9560 7492
rect 8760 5416 9560 6216
rect 8760 -880 9560 -80
rect 7970 -2224 8370 -1824
rect 4370 -3234 4570 -3034
rect -3152 -4577 -2352 -4571
rect -3152 -5377 -3146 -4577
rect -3146 -5377 -2352 -4577
rect -3152 -5383 -2352 -5377
rect 30770 -6490 31170 -6090
rect 31545 -7110 32345 -6510
rect 31540 -7310 32345 -7110
<< metal2 >>
rect 2114 17740 2914 17749
rect 2105 17734 2923 17740
rect 2105 16940 2114 17734
rect 2108 16934 2114 16940
rect 2914 16940 2923 17734
rect 7970 17490 8370 17496
rect 8370 17090 31170 17490
rect 7970 17084 8370 17090
rect 2914 16934 2920 16940
rect 2114 16925 2914 16934
rect 22814 15920 22820 16720
rect 23620 15920 23626 16720
rect 25870 16050 26070 16059
rect -2076 14682 -1276 14691
rect -2076 13873 -1276 13882
rect 8754 11540 8760 12340
rect 9560 11540 9566 12340
rect 8760 10750 9560 10756
rect 22820 10750 23620 15920
rect 30770 15950 31170 17090
rect 9560 9950 10510 10750
rect 22810 9950 24410 10750
rect 8760 9944 9560 9950
rect 8760 8752 9560 8761
rect 7664 7952 8760 8752
rect 8760 7943 9560 7952
rect 8760 7492 9560 7498
rect 7660 6692 8760 7492
rect 8760 6686 9560 6692
rect 25870 6270 26070 15850
rect 29860 15840 31170 15950
rect 29860 15780 31190 15840
rect 29860 15550 31170 15780
rect 8760 6216 9560 6222
rect 7670 5416 8760 6216
rect 24190 6070 26070 6270
rect 8760 5410 9560 5416
rect 7670 4126 8760 4926
rect 9560 4126 9569 4926
rect -1276 3692 -476 3701
rect -3150 3110 -2350 3119
rect -1285 2902 -1276 3692
rect -476 2902 -467 3692
rect 9710 3580 9910 5380
rect 9140 3380 9910 3580
rect 30770 3550 31170 15550
rect -1276 2883 -476 2892
rect 18 2510 24 2696
rect -2350 2496 24 2510
rect 224 2510 230 2696
rect 9140 2510 9340 3380
rect 224 2496 9340 2510
rect -2350 2310 9340 2496
rect 9550 2940 9910 3140
rect -3150 2301 -2350 2310
rect 9550 2100 9750 2940
rect -1640 1900 9750 2100
rect -1640 1690 -1440 1900
rect -2460 1490 -1440 1690
rect -1220 1686 -1020 1695
rect -2460 120 -2260 1490
rect -1220 1477 -1020 1486
rect -2070 1296 -1870 1305
rect -2070 1087 -1870 1096
rect -3159 -680 -3150 120
rect -2350 -680 -2260 120
rect 27640 100 27980 300
rect 8760 -80 9560 -74
rect 9560 -880 10510 -80
rect 8760 -886 9560 -880
rect -502 -1544 -493 -1138
rect -87 -1544 -78 -1138
rect 8765 -1650 9555 -1646
rect 8760 -1655 10060 -1650
rect -2070 -1825 -1870 -1820
rect -1220 -1825 -1020 -1820
rect 7970 -1824 8370 -1818
rect -2074 -2015 -2065 -1825
rect -1875 -2015 -1866 -1825
rect -1224 -2015 -1215 -1825
rect -1025 -2015 -1016 -1825
rect -2070 -4250 -1870 -2015
rect -1220 -4240 -1020 -2015
rect 4170 -2224 7970 -1824
rect 7970 -2230 8370 -2224
rect 4790 -2414 5190 -2408
rect 4170 -2814 4790 -2414
rect 8760 -2445 8765 -1655
rect 9555 -2445 10060 -1655
rect 8760 -2450 10060 -2445
rect 8765 -2454 10060 -2450
rect 4790 -2820 5190 -2814
rect 4370 -3034 4570 -3028
rect 4370 -3240 4570 -3234
rect -499 -3914 -490 -3514
rect -90 -3914 -81 -3514
rect -1220 -4449 -1020 -4440
rect -2070 -4459 -1870 -4450
rect -3152 -4571 -2352 -4565
rect -3161 -5383 -3152 -4571
rect -2352 -5383 -2343 -4571
rect -3152 -5389 -2352 -5383
rect 9260 -6150 10060 -2454
rect 23620 -6150 24420 -4380
rect 27640 -4510 27840 100
rect 27640 -4719 27840 -4710
rect 9260 -6950 24420 -6150
rect 30770 -6090 31170 -3150
rect 30770 -6496 31170 -6490
rect 31540 -6501 31740 300
rect 31540 -6510 32340 -6501
rect 31531 -7310 31540 -6510
rect 32345 -7310 32351 -6510
rect 31550 -7319 32340 -7310
<< via2 >>
rect 2114 16934 2914 17734
rect -2076 13882 -1276 14682
rect 8765 11545 9555 12335
rect 25870 15850 26070 16050
rect 8760 7952 9560 8752
rect 8760 4126 9560 4926
rect -3150 2310 -2350 3110
rect -1276 2892 -476 3692
rect -1220 1486 -1020 1686
rect -2070 1096 -1870 1296
rect -3150 -680 -2350 120
rect -493 -1544 -87 -1138
rect -2065 -2015 -1875 -1825
rect -1215 -2015 -1025 -1825
rect -2070 -4450 -1870 -4250
rect 8765 -2445 9555 -1655
rect -490 -3914 -90 -3514
rect -1220 -4440 -1020 -4240
rect -3152 -5383 -2352 -4571
rect 27640 -4710 27840 -4510
rect 31540 -7110 31545 -6510
rect 31545 -7110 32340 -6510
rect 31540 -7310 32340 -7110
<< metal3 >>
rect 2109 17734 2919 17745
rect 2109 16934 2114 17734
rect 2914 16934 2919 17734
rect 2109 16929 2919 16934
rect 25865 16050 26075 16055
rect 25865 16045 25870 16050
rect 26070 16045 26075 16050
rect 25865 15839 26075 15845
rect -2081 14682 -1271 14687
rect -3150 13882 -2076 14682
rect -1276 13882 -1271 14682
rect -2081 13877 -1271 13882
rect 8760 12335 9560 12340
rect 8760 11545 8765 12335
rect 9555 11545 9560 12335
rect -3150 8180 -476 8980
rect 8760 8757 9560 11545
rect -1276 3697 -476 8180
rect 8755 8752 9565 8757
rect 8755 7952 8760 8752
rect 9560 7952 9565 8752
rect 8755 7947 9565 7952
rect 8755 4926 9565 4931
rect 8755 4126 8760 4926
rect 9560 4126 9565 4926
rect 8755 4121 9565 4126
rect -1281 3692 -471 3697
rect -3155 3110 -2345 3115
rect -3155 2310 -3150 3110
rect -2350 2310 -2345 3110
rect -1281 2892 -1276 3692
rect -476 2892 -471 3692
rect -1281 2887 -471 2892
rect -3155 2305 -2345 2310
rect -1225 1686 -1015 1691
rect -1225 1486 -1220 1686
rect -1020 1486 -1015 1686
rect -1225 1481 -1015 1486
rect -2075 1296 -1865 1301
rect -2075 1096 -2070 1296
rect -1870 1096 -1865 1296
rect -2075 1091 -1865 1096
rect -3155 120 -2345 125
rect -3155 -680 -3150 120
rect -2350 -680 -2345 120
rect -3155 -685 -2345 -680
rect -2070 -1825 -1870 1091
rect -2070 -2015 -2065 -1825
rect -1875 -2015 -1870 -1825
rect -2070 -2020 -1870 -2015
rect -1220 -1825 -1020 1481
rect -498 -1138 -82 -1133
rect -498 -1544 -493 -1138
rect -87 -1544 -82 -1138
rect -498 -1549 -82 -1544
rect -1220 -2015 -1215 -1825
rect -1025 -2015 -1020 -1825
rect -1220 -2020 -1020 -2015
rect -3150 -2307 -2350 -2110
rect -493 -2307 -87 -1549
rect -3150 -2713 -87 -2307
rect 8760 -1655 9560 4121
rect 8760 -2445 8765 -1655
rect 9555 -2445 9560 -1655
rect 8760 -2450 9560 -2445
rect -3150 -2910 -2350 -2713
rect -3150 -3514 -2350 -3310
rect -495 -3514 -85 -3509
rect -3150 -3914 -490 -3514
rect -90 -3914 -85 -3514
rect -3150 -4110 -2350 -3914
rect -495 -3919 -85 -3914
rect -1225 -4240 -1015 -4235
rect -2075 -4250 -1865 -4245
rect -2075 -4450 -2070 -4250
rect -1870 -4450 -1865 -4250
rect -1225 -4440 -1220 -4240
rect -1020 -4440 -160 -4240
rect -1225 -4445 -1015 -4440
rect -2075 -4455 -1865 -4450
rect -3157 -4570 -2347 -4566
rect -3160 -4571 -2347 -4570
rect -3160 -5380 -3152 -4571
rect -3157 -5383 -3152 -5380
rect -2352 -5383 -2347 -4571
rect -3157 -5388 -2347 -5383
rect -2070 -6520 -1870 -4455
rect -360 -6520 -160 -4440
rect 27635 -4505 27845 -4499
rect 27635 -4710 27640 -4705
rect 27840 -4710 27845 -4705
rect 27635 -4715 27845 -4710
rect 31535 -6510 32345 -6505
rect -2370 -7320 -1570 -6520
rect -660 -7320 140 -6520
rect 31535 -7310 31540 -6510
rect 32340 -7310 32345 -6510
rect 31535 -7315 32345 -7310
<< via3 >>
rect 25865 15850 25870 16045
rect 25870 15850 26070 16045
rect 26070 15850 26075 16045
rect 25865 15845 26075 15850
rect 27635 -4510 27845 -4505
rect 27635 -4705 27640 -4510
rect 27640 -4705 27840 -4510
rect 27840 -4705 27845 -4510
<< metal4 >>
rect 25864 16045 26076 16046
rect 25864 15845 25865 16045
rect 26075 15845 26076 16045
rect 25864 15844 26076 15845
rect 25870 -4260 26070 15844
rect 27640 -4504 27840 15660
rect 27634 -4505 27846 -4504
rect 27634 -4705 27635 -4505
rect 27845 -4705 27846 -4505
rect 27634 -4706 27846 -4705
use power_gating  power_gating_0
timestamp 1713815889
transform 1 0 1870 0 1 10256
box -3950 -15173 6766 6365
use schmitt_trigger_pullmid  schmitt_trigger_pullmid_0
timestamp 1713815889
transform 1 0 26390 0 1 -720
box 1390 -3990 5350 16820
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  sky130_fd_pr__cap_mim_m3_1_MPZGNS_0
timestamp 1713813547
transform 1 0 26106 0 1 5700
box -1686 -9960 1686 9960
use vittoz_pierce_osc  vittoz_pierce_osc_0
timestamp 1713815889
transform 1 0 10050 0 1 -2190
box -340 -3540 14370 18841
<< labels >>
flabel metal3 -3150 2310 -2350 3110 0 FreeSans 256 0 0 0 XIN
port 2 nsew
flabel metal3 -3150 -680 -2350 120 0 FreeSans 256 0 0 0 XOUT
port 1 nsew
flabel metal3 -3150 -2914 -2350 -2114 0 FreeSans 256 0 0 0 DVDD
port 7 nsew
flabel metal3 -3150 -4110 -2350 -3310 0 FreeSans 256 0 0 0 DVSS
port 9 nsew
flabel metal3 -3150 8180 -2350 8980 0 FreeSans 256 0 0 0 AVSS
port 8 nsew
flabel metal3 -3150 13881 -2350 14681 0 FreeSans 256 0 0 0 AVDD
port 6 nsew
flabel metal3 2114 16934 2914 17734 0 FreeSans 256 0 0 0 IBIAS
port 10 nsew
flabel metal3 -660 -7320 140 -6520 0 FreeSans 256 0 0 0 STDBY
port 4 nsew
flabel metal3 31540 -7310 32340 -6510 0 FreeSans 256 0 0 0 DOUT
port 5 nsew
flabel metal3 -2370 -7320 -1570 -6520 0 FreeSans 256 0 0 0 ENA
port 3 nsew
flabel metal3 -3162 -5381 -2362 -4581 0 FreeSans 256 0 0 0 GUARD
port 11 nsew
<< end >>
