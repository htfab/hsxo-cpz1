magic
tech sky130A
magscale 1 2
timestamp 1713747467
<< pwell >>
rect -255 -1352 255 1352
<< mvpsubdiff >>
rect -189 1274 189 1286
rect -189 1240 -81 1274
rect 81 1240 189 1274
rect -189 1228 189 1240
rect -189 1178 -131 1228
rect -189 -1178 -177 1178
rect -143 -1178 -131 1178
rect 131 1178 189 1228
rect -189 -1228 -131 -1178
rect 131 -1178 143 1178
rect 177 -1178 189 1178
rect 131 -1228 189 -1178
rect -189 -1240 189 -1228
rect -189 -1274 -81 -1240
rect 81 -1274 189 -1240
rect -189 -1286 189 -1274
<< mvpsubdiffcont >>
rect -81 1240 81 1274
rect -177 -1178 -143 1178
rect 143 -1178 177 1178
rect -81 -1274 81 -1240
<< xpolycontact >>
rect -35 700 35 1132
rect -35 -1132 35 -700
<< xpolyres >>
rect -35 -700 35 700
<< locali >>
rect -177 1240 -81 1274
rect 81 1240 177 1274
rect -177 1178 -143 1240
rect 143 1178 177 1240
rect -177 -1240 -143 -1178
rect 143 -1240 177 -1178
rect -177 -1274 -81 -1240
rect 81 -1274 177 -1240
<< viali >>
rect -19 717 19 1114
rect -19 -1114 19 -717
<< metal1 >>
rect -25 1114 25 1126
rect -25 717 -19 1114
rect 19 717 25 1114
rect -25 705 25 717
rect -25 -717 25 -705
rect -25 -1114 -19 -717
rect 19 -1114 25 -717
rect -25 -1126 25 -1114
<< properties >>
string FIXED_BBOX -160 -1257 160 1257
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 7.16 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 41.989k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
