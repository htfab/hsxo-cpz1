magic
tech sky130A
magscale 1 2
timestamp 1713813547
<< nwell >>
rect 490 2610 5770 2620
rect 490 1830 1120 2610
rect 490 -470 1150 1830
rect 2340 1820 4540 2610
rect 5760 1820 5770 2610
rect 490 -1860 6660 -470
rect 490 -3270 6662 -1860
<< pwell >>
rect 1700 1050 1760 1770
rect 2320 1050 4560 1770
rect 5130 1050 5180 1770
rect 5730 1050 7330 1770
rect 1150 -470 7330 1050
rect 6672 -3270 7330 -470
rect 6040 -6200 7330 -3270
rect 2660 -6830 2810 -6430
rect 1690 -6960 2810 -6830
rect 1690 -7330 2030 -6960
rect 2370 -7304 2390 -7300
rect 2370 -7324 2392 -7304
rect 2400 -7330 2810 -6960
rect 1690 -7460 2810 -7330
rect 4472 -7510 5010 -6210
rect 6672 -7520 7330 -6200
<< locali >>
rect 1630 2924 1830 2930
rect 1630 2736 1636 2924
rect 1824 2736 1830 2924
rect 1630 2556 1830 2736
rect 5050 2924 5250 2930
rect 5050 2736 5056 2924
rect 5244 2736 5250 2924
rect 5050 2556 5250 2736
rect 1184 2550 2282 2556
rect 4604 2550 5702 2556
rect 1178 2482 2288 2550
rect 1178 1952 1252 2482
rect 1604 2350 1862 2482
rect 1604 1952 1678 2350
rect 1178 1884 1678 1952
rect 1788 1952 1862 2350
rect 2214 1952 2288 2482
rect 1788 1884 2288 1952
rect 4598 2482 5708 2550
rect 4598 1952 4672 2482
rect 5024 2350 5282 2482
rect 5024 1952 5098 2350
rect 4598 1884 5098 1952
rect 5208 1952 5282 2350
rect 5634 1952 5708 2482
rect 5208 1884 5708 1952
rect 1184 1878 1672 1884
rect 1794 1878 2282 1884
rect 4604 1878 5092 1884
rect 5214 1878 5702 1884
rect 1184 1734 1672 1738
rect 1794 1734 2282 1738
rect 1184 1732 2282 1734
rect 4604 1732 5092 1738
rect 5214 1732 5702 1738
rect 1178 1664 2288 1732
rect 1178 1152 1252 1664
rect 1604 1546 1862 1664
rect 1604 1152 1678 1546
rect 1178 1084 1678 1152
rect 1788 1152 1862 1546
rect 2214 1152 2288 1664
rect 1788 1084 2288 1152
rect 4598 1664 5098 1732
rect 4598 1152 4672 1664
rect 5024 1280 5098 1664
rect 5208 1664 5708 1732
rect 5208 1280 5282 1664
rect 5024 1152 5282 1280
rect 5634 1152 5708 1664
rect 4598 1084 5708 1152
rect 1184 1078 1672 1084
rect 1794 1078 2282 1084
rect 4604 1078 5702 1084
rect 5050 774 5250 1078
rect 5050 586 5056 774
rect 5244 586 5250 774
rect 5050 580 5250 586
rect 3260 -1724 3266 -1530
rect 4054 -1724 4060 -1680
rect 3260 -1840 4060 -1724
rect 3260 -1920 4692 -1840
rect 2410 -1924 2882 -1920
rect 3160 -1924 5040 -1920
rect 874 -1930 6598 -1924
rect 868 -1998 6604 -1930
rect 868 -3128 942 -1998
rect 2400 -3128 2902 -1998
rect 4360 -2120 5072 -1998
rect 4360 -3128 4434 -2120
rect 868 -3130 4434 -3128
rect 570 -3196 4434 -3130
rect 4998 -3128 5072 -2120
rect 6530 -3128 6604 -1998
rect 4998 -3196 6604 -3128
rect 570 -3200 4428 -3196
rect 570 -3202 2468 -3200
rect 2834 -3202 4428 -3200
rect 5004 -3202 6598 -3196
rect 570 -3330 1770 -3202
rect 570 -3550 590 -3330
rect 1750 -3550 1770 -3330
rect 570 -3560 1770 -3550
rect 2844 -6238 4438 -6232
rect 5044 -6238 6638 -6232
rect 2838 -6306 4444 -6238
rect 965 -6750 1781 -6739
rect 965 -6830 980 -6750
rect 1060 -6830 1690 -6750
rect 1770 -6830 1781 -6750
rect 965 -6840 1781 -6830
rect 965 -7450 1070 -6840
rect 1175 -6950 1571 -6949
rect 1175 -7040 1290 -6950
rect 1450 -7040 1571 -6950
rect 1175 -7049 1571 -7040
rect 1175 -7245 1275 -7049
rect 1471 -7245 1571 -7049
rect 1175 -7345 1571 -7245
rect 1680 -7450 1781 -6840
rect 2010 -6960 2414 -6945
rect 2010 -7030 2020 -6960
rect 2090 -7030 2330 -6960
rect 2400 -7030 2414 -6960
rect 2010 -7045 2414 -7030
rect 2010 -7249 2112 -7045
rect 2314 -7249 2414 -7045
rect 2010 -7270 2414 -7249
rect 2010 -7340 2020 -7270
rect 2090 -7340 2330 -7270
rect 2400 -7340 2414 -7270
rect 2010 -7349 2414 -7340
rect 965 -7460 1781 -7450
rect 2838 -7418 2912 -6306
rect 4370 -7295 4444 -6306
rect 5038 -6306 6644 -6238
rect 5038 -7295 5112 -6306
rect 4370 -7418 5112 -7295
rect 6570 -7418 6644 -6306
rect 2838 -7460 6644 -7418
rect 965 -7540 980 -7460
rect 1060 -7540 1690 -7460
rect 1770 -7540 1781 -7460
rect 965 -7555 1781 -7540
rect 2320 -7466 6644 -7460
rect 2320 -7654 2326 -7466
rect 2514 -7486 6644 -7466
rect 2514 -7492 6638 -7486
rect 2514 -7654 2890 -7492
rect 4392 -7500 5092 -7492
rect 2320 -7660 2890 -7654
<< viali >>
rect 1636 2736 1824 2924
rect 5056 2736 5244 2924
rect 5056 586 5244 774
rect 3266 -1724 4054 -936
rect 590 -3550 1750 -3330
rect 980 -6830 1060 -6750
rect 1690 -6830 1770 -6750
rect 1290 -7040 1450 -6950
rect 2020 -7030 2090 -6960
rect 2330 -7030 2400 -6960
rect 2020 -7340 2090 -7270
rect 2330 -7340 2400 -7270
rect 980 -7540 1060 -7460
rect 1690 -7540 1770 -7460
rect 2326 -7654 2514 -7466
<< metal1 >>
rect -270 3530 530 3536
rect -276 2730 -270 2930
rect 1630 2930 1830 2936
rect 1624 2730 1630 2930
rect 1830 2730 1836 2930
rect -270 -3320 530 2730
rect 1630 2724 1830 2730
rect 722 1727 728 1932
rect 933 1727 939 1932
rect 2300 1730 2440 1930
rect 2542 1727 2548 1932
rect 2753 1727 2759 1932
rect 728 -1920 933 1727
rect 1934 940 1940 1140
rect 2140 940 2146 1140
rect 1940 780 2140 940
rect 1104 580 1110 780
rect 1310 580 2140 780
rect 2548 -1538 2753 1727
rect 2900 -1160 3100 3936
rect 3254 2730 3260 3530
rect 4060 2730 4066 3530
rect 5050 2930 5250 2936
rect 5044 2730 5050 2930
rect 5250 2730 5256 2930
rect 3260 -930 4060 2730
rect 5050 2724 5250 2730
rect 4318 1930 4503 1932
rect 6542 1930 6742 1936
rect 4318 1730 4360 1930
rect 4560 1730 4590 1930
rect 6537 1730 6542 1902
rect 4318 -928 4523 1730
rect 4744 934 4750 1134
rect 4950 934 4956 1134
rect 5354 940 5360 1140
rect 5560 940 5566 1140
rect 4750 -180 4950 934
rect 5050 780 5250 786
rect 5050 574 5250 580
rect 4750 -386 4950 -380
rect 5360 -540 5560 940
rect 5360 -746 5560 -740
rect 2894 -1360 2900 -1160
rect 3100 -1360 3106 -1160
rect 2542 -1743 2548 -1538
rect 2753 -1743 2759 -1538
rect 4312 -1133 4318 -928
rect 4523 -1133 4529 -928
rect 3260 -1736 4060 -1730
rect 6537 -1920 6742 1730
rect 7350 780 8150 3536
rect 7344 -20 7350 780
rect 8150 -20 8156 780
rect 6969 -928 7174 -922
rect 6961 -1133 6967 -928
rect 7172 -1133 7178 -928
rect 6967 -1362 7174 -1133
rect 728 -2122 4572 -1920
rect 730 -2125 4572 -2122
rect 730 -3005 935 -2125
rect 1012 -2175 1066 -2165
rect 1012 -2329 1066 -2319
rect 1328 -2175 1382 -2165
rect 1328 -2329 1382 -2319
rect 1644 -2175 1698 -2165
rect 1644 -2329 1698 -2319
rect 1960 -2175 2014 -2165
rect 1960 -2329 2014 -2319
rect 2276 -2175 2330 -2165
rect 2276 -2329 2330 -2319
rect 1170 -2807 1224 -2797
rect 1170 -2961 1224 -2951
rect 1486 -2807 1540 -2797
rect 1486 -2961 1540 -2951
rect 1802 -2807 1856 -2797
rect 1802 -2961 1856 -2951
rect 2118 -2807 2172 -2797
rect 2118 -2961 2172 -2951
rect 2407 -3005 2895 -2125
rect 2972 -2175 3026 -2165
rect 2972 -2329 3026 -2319
rect 3288 -2175 3342 -2165
rect 3288 -2329 3342 -2319
rect 3604 -2175 3658 -2165
rect 3604 -2329 3658 -2319
rect 3920 -2175 3974 -2165
rect 3920 -2329 3974 -2319
rect 4236 -2175 4290 -2165
rect 4236 -2329 4290 -2319
rect 3130 -2807 3184 -2797
rect 3130 -2961 3184 -2951
rect 3446 -2807 3500 -2797
rect 3446 -2961 3500 -2951
rect 3762 -2807 3816 -2797
rect 3762 -2961 3816 -2951
rect 4078 -2807 4132 -2797
rect 4078 -2961 4132 -2951
rect 4367 -3005 4572 -2125
rect 730 -3210 4572 -3005
rect 4860 -2125 6742 -1920
rect 4860 -3005 5065 -2125
rect 5142 -2175 5196 -2165
rect 5142 -2329 5196 -2319
rect 5458 -2175 5512 -2165
rect 5458 -2329 5512 -2319
rect 5774 -2175 5828 -2165
rect 5774 -2329 5828 -2319
rect 6090 -2175 6144 -2165
rect 6090 -2329 6144 -2319
rect 6406 -2175 6460 -2165
rect 6406 -2329 6460 -2319
rect 5300 -2807 5354 -2797
rect 5300 -2961 5354 -2951
rect 5616 -2807 5670 -2797
rect 5616 -2961 5670 -2951
rect 5932 -2807 5986 -2797
rect 5932 -2961 5986 -2951
rect 6248 -2807 6302 -2797
rect 6248 -2961 6302 -2951
rect 6537 -3005 6742 -2125
rect 4860 -3210 6742 -3005
rect -270 -3330 1770 -3320
rect -270 -3550 590 -3330
rect 1750 -3550 1770 -3330
rect -270 -4120 1770 -3550
rect 970 -6510 1770 -4120
rect 2542 -6303 2548 -6098
rect 2753 -6220 2895 -6098
rect 6969 -6220 7174 -1362
rect 2753 -6303 4572 -6220
rect 2690 -6425 4572 -6303
rect 915 -6750 1115 -6700
rect 915 -6830 980 -6750
rect 1060 -6830 1115 -6750
rect 510 -7050 710 -7044
rect -1586 -7250 -1580 -7050
rect -1380 -7250 -1374 -7050
rect -1156 -7250 -1150 -7050
rect -950 -7250 -944 -7050
rect -736 -7250 -730 -7050
rect -530 -7250 -524 -7050
rect -316 -7250 -310 -7050
rect -110 -7250 -104 -7050
rect 84 -7250 90 -7050
rect 290 -7250 296 -7050
rect 710 -7250 716 -7050
rect -1580 -8666 -1380 -7250
rect -1150 -8666 -950 -7250
rect -730 -8666 -530 -7250
rect -310 -8666 -110 -7250
rect 90 -8666 290 -7250
rect 510 -8656 710 -7250
rect 915 -7405 1115 -6830
rect 1271 -6950 1471 -6510
rect 1271 -7040 1290 -6950
rect 1450 -7040 1471 -6950
rect 1271 -7050 1471 -7040
rect 1631 -6750 1831 -6690
rect 1631 -6830 1690 -6750
rect 1770 -6830 1831 -6750
rect 1300 -7090 1440 -7080
rect 1300 -7210 1310 -7090
rect 1430 -7210 1440 -7090
rect 1300 -7220 1440 -7210
rect 1631 -7260 1831 -6830
rect 1900 -6960 2520 -6840
rect 1900 -7030 2020 -6960
rect 2090 -7030 2330 -6960
rect 2400 -7030 2520 -6960
rect 1900 -7040 2520 -7030
rect 1900 -7260 2100 -7040
rect 2140 -7090 2280 -7080
rect 2140 -7210 2150 -7090
rect 2270 -7210 2280 -7090
rect 2140 -7220 2280 -7210
rect 2320 -7260 2520 -7040
rect 1631 -7270 2520 -7260
rect 1631 -7340 2020 -7270
rect 2090 -7340 2330 -7270
rect 2400 -7340 2520 -7270
rect 1631 -7405 2520 -7340
rect 915 -7460 2520 -7405
rect 2690 -7295 2890 -6425
rect 2982 -6474 3036 -6464
rect 2982 -6628 3036 -6618
rect 3298 -6474 3352 -6464
rect 3298 -6628 3352 -6618
rect 3614 -6474 3668 -6464
rect 3614 -6628 3668 -6618
rect 3930 -6474 3984 -6464
rect 3930 -6628 3984 -6618
rect 4246 -6474 4300 -6464
rect 4246 -6628 4300 -6618
rect 3140 -7106 3194 -7096
rect 3140 -7260 3194 -7250
rect 3456 -7106 3510 -7096
rect 3456 -7260 3510 -7250
rect 3772 -7106 3826 -7096
rect 3772 -7260 3826 -7250
rect 4088 -7106 4142 -7096
rect 4088 -7260 4142 -7250
rect 4372 -7295 4572 -6425
rect 915 -7605 954 -7460
rect 1154 -7540 1690 -7460
rect 1770 -7540 1831 -7460
rect 948 -7660 954 -7605
rect 1154 -7605 1831 -7540
rect 1154 -7660 1160 -7605
rect 2314 -7660 2320 -7460
rect 2520 -7660 2526 -7460
rect 2690 -7500 4572 -7295
rect 4870 -6425 7174 -6220
rect 4870 -7295 5070 -6425
rect 5182 -6474 5236 -6464
rect 5182 -6628 5236 -6618
rect 5498 -6474 5552 -6464
rect 5498 -6628 5552 -6618
rect 5814 -6474 5868 -6464
rect 5814 -6628 5868 -6618
rect 6130 -6474 6184 -6464
rect 6130 -6628 6184 -6618
rect 6446 -6474 6500 -6464
rect 6446 -6628 6500 -6618
rect 5340 -7106 5394 -7096
rect 5340 -7260 5394 -7250
rect 5656 -7106 5710 -7096
rect 5656 -7260 5710 -7250
rect 5972 -7106 6026 -7096
rect 5972 -7260 6026 -7250
rect 6288 -7106 6342 -7096
rect 6288 -7260 6342 -7250
rect 6532 -7295 6732 -6425
rect 7350 -7290 8150 -20
rect 4870 -7500 6732 -7295
rect 2320 -7666 2520 -7660
rect 7344 -8090 7350 -7290
rect 8150 -8090 8156 -7290
rect 7350 -8096 8150 -8090
<< via1 >>
rect -270 2730 530 3530
rect 1630 2924 1830 2930
rect 1630 2736 1636 2924
rect 1636 2736 1824 2924
rect 1824 2736 1830 2924
rect 1630 2730 1830 2736
rect 728 1727 933 1932
rect 2548 1727 2753 1932
rect 1940 940 2140 1140
rect 1110 580 1310 780
rect 3260 2730 4060 3530
rect 5050 2924 5250 2930
rect 5050 2736 5056 2924
rect 5056 2736 5244 2924
rect 5244 2736 5250 2924
rect 5050 2730 5250 2736
rect 4360 1730 4560 1930
rect 6542 1730 6742 1930
rect 4750 934 4950 1134
rect 5360 940 5560 1140
rect 5050 774 5250 780
rect 5050 586 5056 774
rect 5056 586 5244 774
rect 5244 586 5250 774
rect 5050 580 5250 586
rect 4750 -380 4950 -180
rect 5360 -740 5560 -540
rect 3260 -936 4060 -930
rect 2900 -1360 3100 -1160
rect 2548 -1743 2753 -1538
rect 3260 -1724 3266 -936
rect 3266 -1724 4054 -936
rect 4054 -1724 4060 -936
rect 4318 -1133 4523 -928
rect 3260 -1730 4060 -1724
rect 7350 -20 8150 780
rect 6967 -1133 7172 -928
rect 1012 -2319 1066 -2175
rect 1328 -2319 1382 -2175
rect 1644 -2319 1698 -2175
rect 1960 -2319 2014 -2175
rect 2276 -2319 2330 -2175
rect 1170 -2951 1224 -2807
rect 1486 -2951 1540 -2807
rect 1802 -2951 1856 -2807
rect 2118 -2951 2172 -2807
rect 2972 -2319 3026 -2175
rect 3288 -2319 3342 -2175
rect 3604 -2319 3658 -2175
rect 3920 -2319 3974 -2175
rect 4236 -2319 4290 -2175
rect 3130 -2951 3184 -2807
rect 3446 -2951 3500 -2807
rect 3762 -2951 3816 -2807
rect 4078 -2951 4132 -2807
rect 5142 -2319 5196 -2175
rect 5458 -2319 5512 -2175
rect 5774 -2319 5828 -2175
rect 6090 -2319 6144 -2175
rect 6406 -2319 6460 -2175
rect 5300 -2951 5354 -2807
rect 5616 -2951 5670 -2807
rect 5932 -2951 5986 -2807
rect 6248 -2951 6302 -2807
rect 2548 -6303 2753 -6098
rect -1580 -7250 -1380 -7050
rect -1150 -7250 -950 -7050
rect -730 -7250 -530 -7050
rect -310 -7250 -110 -7050
rect 90 -7250 290 -7050
rect 510 -7250 710 -7050
rect 1310 -7210 1430 -7090
rect 2150 -7210 2270 -7090
rect 2982 -6618 3036 -6474
rect 3298 -6618 3352 -6474
rect 3614 -6618 3668 -6474
rect 3930 -6618 3984 -6474
rect 4246 -6618 4300 -6474
rect 3140 -7250 3194 -7106
rect 3456 -7250 3510 -7106
rect 3772 -7250 3826 -7106
rect 4088 -7250 4142 -7106
rect 954 -7540 980 -7460
rect 980 -7540 1060 -7460
rect 1060 -7540 1154 -7460
rect 954 -7660 1154 -7540
rect 2320 -7466 2520 -7460
rect 2320 -7654 2326 -7466
rect 2326 -7654 2514 -7466
rect 2514 -7654 2520 -7466
rect 2320 -7660 2520 -7654
rect 5182 -6618 5236 -6474
rect 5498 -6618 5552 -6474
rect 5814 -6618 5868 -6474
rect 6130 -6618 6184 -6474
rect 6446 -6618 6500 -6474
rect 5340 -7250 5394 -7106
rect 5656 -7250 5710 -7106
rect 5972 -7250 6026 -7106
rect 6288 -7250 6342 -7106
rect 7350 -8090 8150 -7290
<< metal2 >>
rect 3260 3530 4060 3536
rect -1590 3525 -270 3530
rect -1594 2735 -270 3525
rect -1590 2730 -270 2735
rect 530 2930 3260 3530
rect 530 2730 1630 2930
rect 1830 2730 3260 2930
rect 4060 2930 5850 3530
rect 4060 2730 5050 2930
rect 5250 2730 5850 2930
rect -270 2724 -70 2730
rect 1630 2500 1830 2730
rect 3260 2724 4060 2730
rect 5050 2500 5250 2730
rect 728 1932 933 1938
rect 2548 1932 2753 1938
rect 933 1727 1172 1932
rect 2388 1930 2548 1932
rect 2250 1730 2548 1930
rect 2388 1727 2548 1730
rect 728 1721 933 1727
rect 2548 1721 2753 1727
rect 4360 1930 4560 1936
rect 4560 1730 4640 1930
rect 5670 1730 6542 1930
rect 6742 1730 6748 1930
rect 4360 1724 4560 1730
rect 1940 1140 2140 1146
rect -1580 940 1530 1140
rect -1580 -7050 -1380 940
rect 1110 780 1310 786
rect -1580 -7256 -1380 -7250
rect -1150 580 1110 780
rect -1150 -7050 -950 580
rect 1110 574 1310 580
rect 1630 780 1830 1120
rect 1940 934 2140 940
rect 4750 1134 4950 1146
rect 5360 1140 5560 1146
rect 4750 928 4950 934
rect 5050 780 5250 1140
rect 5360 934 5560 940
rect 7350 780 8150 786
rect 1630 580 5050 780
rect 5250 580 7350 780
rect 1630 -20 7350 580
rect 7350 -26 8150 -20
rect -1150 -7256 -950 -7250
rect -730 -380 4750 -180
rect 4950 -380 4956 -180
rect -730 -7050 -530 -380
rect -730 -7256 -530 -7250
rect -310 -740 5360 -540
rect 5560 -740 5566 -540
rect -310 -7050 -110 -740
rect 4318 -928 4523 -922
rect 6967 -928 7172 -922
rect 2900 -1160 3100 -1154
rect 2140 -1360 2900 -1160
rect 2140 -2130 2340 -1360
rect 2900 -1366 3100 -1360
rect 3254 -1510 3260 -930
rect 2548 -1538 2753 -1532
rect 4060 -1530 4066 -930
rect 4523 -1133 6967 -928
rect 7172 -1133 7180 -928
rect 4318 -1139 4523 -1133
rect 6967 -1139 7172 -1133
rect 4060 -1730 6472 -1530
rect 1000 -2175 2342 -2130
rect 1000 -2319 1012 -2175
rect 1066 -2319 1328 -2175
rect 1382 -2319 1644 -2175
rect 1698 -2319 1960 -2175
rect 2014 -2319 2276 -2175
rect 2330 -2319 2342 -2175
rect 1000 -2330 2342 -2319
rect -310 -7256 -110 -7250
rect 90 -2807 2342 -2800
rect 90 -2951 1170 -2807
rect 1224 -2951 1486 -2807
rect 1540 -2951 1802 -2807
rect 1856 -2951 2118 -2807
rect 2172 -2951 2342 -2807
rect 90 -3000 2342 -2951
rect 90 -7050 290 -3000
rect 2548 -6098 2753 -1743
rect 2960 -2175 6472 -1730
rect 2960 -2319 2972 -2175
rect 3026 -2319 3288 -2175
rect 3342 -2319 3604 -2175
rect 3658 -2319 3920 -2175
rect 3974 -2319 4236 -2175
rect 4290 -2319 5142 -2175
rect 5196 -2319 5458 -2175
rect 5512 -2319 5774 -2175
rect 5828 -2319 6090 -2175
rect 6144 -2319 6406 -2175
rect 6460 -2319 6472 -2175
rect 2960 -2330 6472 -2319
rect 6700 -2800 8950 -2400
rect 2960 -2807 4392 -2800
rect 2960 -2951 3130 -2807
rect 3184 -2951 3446 -2807
rect 3500 -2951 3762 -2807
rect 3816 -2951 4078 -2807
rect 4132 -2951 4392 -2807
rect 2960 -3450 4392 -2951
rect 5130 -2807 8950 -2800
rect 5130 -2951 5300 -2807
rect 5354 -2951 5616 -2807
rect 5670 -2951 5932 -2807
rect 5986 -2951 6248 -2807
rect 6302 -2951 8950 -2807
rect 5130 -3200 8950 -2951
rect 5130 -3300 7500 -3200
rect 3590 -3660 4392 -3450
rect 3590 -4460 8950 -3660
rect 3580 -5740 8950 -4940
rect 3580 -6160 4380 -5740
rect 2548 -6309 2753 -6303
rect 2970 -6474 4402 -6160
rect 2970 -6618 2982 -6474
rect 3036 -6618 3298 -6474
rect 3352 -6618 3614 -6474
rect 3668 -6618 3930 -6474
rect 3984 -6618 4246 -6474
rect 4300 -6618 4402 -6474
rect 2970 -6630 4402 -6618
rect 5170 -6230 7500 -6150
rect 5170 -6474 8950 -6230
rect 5170 -6618 5182 -6474
rect 5236 -6618 5498 -6474
rect 5552 -6618 5814 -6474
rect 5868 -6618 6130 -6474
rect 6184 -6618 6446 -6474
rect 6500 -6618 8950 -6474
rect 5170 -6630 8950 -6618
rect 6700 -7030 8950 -6630
rect 510 -7050 710 -7044
rect 1271 -7050 1471 -7049
rect 504 -7250 510 -7050
rect 710 -7090 2310 -7050
rect 710 -7210 1310 -7090
rect 1430 -7210 2150 -7090
rect 2270 -7210 2310 -7090
rect 710 -7250 2310 -7210
rect 2970 -7106 6522 -7100
rect 2970 -7250 3140 -7106
rect 3194 -7250 3456 -7106
rect 3510 -7250 3772 -7106
rect 3826 -7250 4088 -7106
rect 4142 -7250 5340 -7106
rect 5394 -7250 5656 -7106
rect 5710 -7250 5972 -7106
rect 6026 -7250 6288 -7106
rect 6342 -7250 6522 -7106
rect 90 -7256 290 -7250
rect 510 -7256 710 -7250
rect 2970 -7290 6522 -7250
rect 7350 -7290 8150 -7284
rect 954 -7460 1154 -7454
rect 2320 -7460 2520 -7454
rect 2970 -7460 7350 -7290
rect -790 -7660 954 -7460
rect 1154 -7660 2320 -7460
rect 2520 -7660 7350 -7460
rect -790 -8090 7350 -7660
rect 8150 -8090 8156 -7290
rect -790 -8260 3770 -8090
rect 7350 -8096 8150 -8090
use level_shifter_ad  level_shifter_ad_0
timestamp 1713804741
transform 1 0 140 0 1 2910
box 880 -1970 2310 -210
use level_shifter_ad  level_shifter_ad_1
timestamp 1713804741
transform 1 0 3560 0 1 2910
box 880 -1970 2310 -210
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_0
timestamp 1713804741
transform 1 0 1373 0 1 -7147
box -423 -423 423 423
use sky130_fd_pr__diode_pw2nd_11v0_FT76RJ  sky130_fd_pr__diode_pw2nd_11v0_FT76RJ_0
timestamp 1713804741
transform 1 0 2212 0 1 -7147
box -217 -217 217 217
use sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ  sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ_0
timestamp 1713804741
transform 1 0 3641 0 1 -6862
box -831 -658 831 658
use sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ  sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ_1
timestamp 1713804741
transform 1 0 5841 0 1 -6862
box -831 -658 831 658
use sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6  sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6_0
timestamp 1713804741
transform 1 0 1671 0 1 -2563
box -861 -697 861 697
use sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6  XM1
timestamp 1713804741
transform 1 0 5801 0 1 -2563
box -861 -697 861 697
use sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6  XM25
timestamp 1713804741
transform 1 0 3631 0 1 -2563
box -861 -697 861 697
<< labels >>
flabel metal2 8150 -5740 8950 -4940 0 FreeSans 256 0 0 0 EG_AVSS
port 7 nsew
flabel metal2 8150 -3200 8950 -2400 0 FreeSans 256 0 0 0 SG_AVDD
port 8 nsew
flabel metal1 7350 2730 8150 3530 0 FreeSans 256 0 0 0 AVSS
port 2 nsew
flabel metal2 8150 -4460 8950 -3660 0 FreeSans 256 0 0 0 EG_AVDD
port 6 nsew
flabel metal2 8150 -7030 8950 -6230 0 FreeSans 256 0 0 0 SG_AVSS
port 9 nsew
flabel metal1 2900 3730 3100 3930 0 FreeSans 256 0 0 0 IBIAS
port 5 nsew
flabel metal1 510 -8650 710 -8450 0 FreeSans 256 0 0 0 XIN
port 11 nsew
flabel metal1 90 -8660 290 -8460 0 FreeSans 256 0 0 0 EG_IBIAS
port 10 nsew
flabel metal1 -310 -8660 -110 -8460 0 FreeSans 256 0 0 0 STDBY_B
port 13 nsew
flabel metal1 -1150 -8660 -950 -8460 0 FreeSans 256 0 0 0 ENA_B
port 12 nsew
flabel metal1 -730 -8660 -530 -8460 0 FreeSans 256 0 0 0 STDBY
port 4 nsew
flabel metal1 -1580 -8660 -1380 -8460 0 FreeSans 256 0 0 0 ENA
port 3 nsew
flabel metal2 -1590 2730 -790 3530 0 FreeSans 256 0 0 0 AVDD
port 1 nsew
flabel metal2 5050 2730 5850 3530 0 FreeSans 256 0 0 0 AVDD
port 1 nsew
flabel metal2 -790 -8260 10 -7460 0 FreeSans 256 0 0 0 AVSS
port 2 nsew
<< end >>
