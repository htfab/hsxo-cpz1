magic
tech sky130A
magscale 1 2
timestamp 1713784524
<< nwell >>
rect -861 -697 861 697
<< mvpmos >>
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
<< mvpdiff >>
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
<< mvpdiffc >>
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
<< mvnsubdiff >>
rect -795 619 795 631
rect -795 585 -687 619
rect 687 585 795 619
rect -795 573 795 585
rect -795 523 -737 573
rect -795 -523 -783 523
rect -749 -523 -737 523
rect 737 523 795 573
rect -795 -573 -737 -523
rect 737 -523 749 523
rect 783 -523 795 523
rect 737 -573 795 -523
rect -795 -585 795 -573
rect -795 -619 -687 -585
rect 687 -619 795 -585
rect -795 -631 795 -619
<< mvnsubdiffcont >>
rect -687 585 687 619
rect -783 -523 -749 523
rect 749 -523 783 523
rect -687 -619 687 -585
<< poly >>
rect -603 481 -503 497
rect -603 447 -587 481
rect -519 447 -503 481
rect -603 400 -503 447
rect -445 481 -345 497
rect -445 447 -429 481
rect -361 447 -345 481
rect -445 400 -345 447
rect -287 481 -187 497
rect -287 447 -271 481
rect -203 447 -187 481
rect -287 400 -187 447
rect -129 481 -29 497
rect -129 447 -113 481
rect -45 447 -29 481
rect -129 400 -29 447
rect 29 481 129 497
rect 29 447 45 481
rect 113 447 129 481
rect 29 400 129 447
rect 187 481 287 497
rect 187 447 203 481
rect 271 447 287 481
rect 187 400 287 447
rect 345 481 445 497
rect 345 447 361 481
rect 429 447 445 481
rect 345 400 445 447
rect 503 481 603 497
rect 503 447 519 481
rect 587 447 603 481
rect 503 400 603 447
rect -603 -447 -503 -400
rect -603 -481 -587 -447
rect -519 -481 -503 -447
rect -603 -497 -503 -481
rect -445 -447 -345 -400
rect -445 -481 -429 -447
rect -361 -481 -345 -447
rect -445 -497 -345 -481
rect -287 -447 -187 -400
rect -287 -481 -271 -447
rect -203 -481 -187 -447
rect -287 -497 -187 -481
rect -129 -447 -29 -400
rect -129 -481 -113 -447
rect -45 -481 -29 -447
rect -129 -497 -29 -481
rect 29 -447 129 -400
rect 29 -481 45 -447
rect 113 -481 129 -447
rect 29 -497 129 -481
rect 187 -447 287 -400
rect 187 -481 203 -447
rect 271 -481 287 -447
rect 187 -497 287 -481
rect 345 -447 445 -400
rect 345 -481 361 -447
rect 429 -481 445 -447
rect 345 -497 445 -481
rect 503 -447 603 -400
rect 503 -481 519 -447
rect 587 -481 603 -447
rect 503 -497 603 -481
<< polycont >>
rect -587 447 -519 481
rect -429 447 -361 481
rect -271 447 -203 481
rect -113 447 -45 481
rect 45 447 113 481
rect 203 447 271 481
rect 361 447 429 481
rect 519 447 587 481
rect -587 -481 -519 -447
rect -429 -481 -361 -447
rect -271 -481 -203 -447
rect -113 -481 -45 -447
rect 45 -481 113 -447
rect 203 -481 271 -447
rect 361 -481 429 -447
rect 519 -481 587 -447
<< locali >>
rect -783 585 -687 619
rect 687 585 783 619
rect -783 523 -749 585
rect 749 523 783 585
rect -603 447 -587 481
rect -519 447 -503 481
rect -445 447 -429 481
rect -361 447 -345 481
rect -287 447 -271 481
rect -203 447 -187 481
rect -129 447 -113 481
rect -45 447 -29 481
rect 29 447 45 481
rect 113 447 129 481
rect 187 447 203 481
rect 271 447 287 481
rect 345 447 361 481
rect 429 447 445 481
rect 503 447 519 481
rect 587 447 603 481
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect -603 -481 -587 -447
rect -519 -481 -503 -447
rect -445 -481 -429 -447
rect -361 -481 -345 -447
rect -287 -481 -271 -447
rect -203 -481 -187 -447
rect -129 -481 -113 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 113 -481 129 -447
rect 187 -481 203 -447
rect 271 -481 287 -447
rect 345 -481 361 -447
rect 429 -481 445 -447
rect 503 -481 519 -447
rect 587 -481 603 -447
rect -783 -585 -749 -523
rect 749 -585 783 -523
rect -783 -619 -687 -585
rect 687 -619 783 -585
<< viali >>
rect -587 447 -519 481
rect -429 447 -361 481
rect -271 447 -203 481
rect -113 447 -45 481
rect 45 447 113 481
rect 203 447 271 481
rect 361 447 429 481
rect 519 447 587 481
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect -587 -481 -519 -447
rect -429 -481 -361 -447
rect -271 -481 -203 -447
rect -113 -481 -45 -447
rect 45 -481 113 -447
rect 203 -481 271 -447
rect 361 -481 429 -447
rect 519 -481 587 -447
<< metal1 >>
rect -599 481 -507 487
rect -599 447 -587 481
rect -519 447 -507 481
rect -599 441 -507 447
rect -441 481 -349 487
rect -441 447 -429 481
rect -361 447 -349 481
rect -441 441 -349 447
rect -283 481 -191 487
rect -283 447 -271 481
rect -203 447 -191 481
rect -283 441 -191 447
rect -125 481 -33 487
rect -125 447 -113 481
rect -45 447 -33 481
rect -125 441 -33 447
rect 33 481 125 487
rect 33 447 45 481
rect 113 447 125 481
rect 33 441 125 447
rect 191 481 283 487
rect 191 447 203 481
rect 271 447 283 481
rect 191 441 283 447
rect 349 481 441 487
rect 349 447 361 481
rect 429 447 441 481
rect 349 441 441 447
rect 507 481 599 487
rect 507 447 519 481
rect 587 447 599 481
rect 507 441 599 447
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect -599 -447 -507 -441
rect -599 -481 -587 -447
rect -519 -481 -507 -447
rect -599 -487 -507 -481
rect -441 -447 -349 -441
rect -441 -481 -429 -447
rect -361 -481 -349 -447
rect -441 -487 -349 -481
rect -283 -447 -191 -441
rect -283 -481 -271 -447
rect -203 -481 -191 -447
rect -283 -487 -191 -481
rect -125 -447 -33 -441
rect -125 -481 -113 -447
rect -45 -481 -33 -447
rect -125 -487 -33 -481
rect 33 -447 125 -441
rect 33 -481 45 -447
rect 113 -481 125 -447
rect 33 -487 125 -481
rect 191 -447 283 -441
rect 191 -481 203 -447
rect 271 -481 283 -447
rect 191 -487 283 -481
rect 349 -447 441 -441
rect 349 -481 361 -447
rect 429 -481 441 -447
rect 349 -487 441 -481
rect 507 -447 599 -441
rect 507 -481 519 -447
rect 587 -481 599 -447
rect 507 -487 599 -481
<< properties >>
string FIXED_BBOX -766 -602 766 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
