magic
tech sky130A
magscale 1 2
timestamp 1713747467
<< pwell >>
rect -255 -932 255 932
<< mvpsubdiff >>
rect -189 854 189 866
rect -189 820 -81 854
rect 81 820 189 854
rect -189 808 189 820
rect -189 758 -131 808
rect -189 -758 -177 758
rect -143 -758 -131 758
rect 131 758 189 808
rect -189 -808 -131 -758
rect 131 -758 143 758
rect 177 -758 189 758
rect 131 -808 189 -758
rect -189 -820 189 -808
rect -189 -854 -81 -820
rect 81 -854 189 -820
rect -189 -866 189 -854
<< mvpsubdiffcont >>
rect -81 820 81 854
rect -177 -758 -143 758
rect 143 -758 177 758
rect -81 -854 81 -820
<< xpolycontact >>
rect -35 280 35 712
rect -35 -712 35 -280
<< xpolyres >>
rect -35 -280 35 280
<< locali >>
rect -177 820 -81 854
rect 81 820 177 854
rect -177 758 -143 820
rect 143 758 177 820
rect -177 -820 -143 -758
rect 143 -820 177 -758
rect -177 -854 -81 -820
rect 81 -854 177 -820
<< viali >>
rect -19 297 19 694
rect -19 -694 19 -297
<< metal1 >>
rect -25 694 25 706
rect -25 297 -19 694
rect 19 297 25 694
rect -25 285 25 297
rect -25 -297 25 -285
rect -25 -694 -19 -297
rect 19 -694 25 -297
rect -25 -706 25 -694
<< properties >>
string FIXED_BBOX -160 -837 160 837
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2.96 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 17.989k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
