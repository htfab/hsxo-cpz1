magic
tech sky130A
magscale 1 2
timestamp 1712821206
<< pwell >>
rect -201 -878 201 878
<< psubdiff >>
rect -165 808 -69 842
rect 69 808 165 842
rect -165 746 -131 808
rect 131 746 165 808
rect -165 -808 -131 -746
rect 131 -808 165 -746
rect -165 -842 -69 -808
rect 69 -842 165 -808
<< psubdiffcont >>
rect -69 808 69 842
rect -165 -746 -131 746
rect 131 -746 165 746
rect -69 -842 69 -808
<< xpolycontact >>
rect -35 280 35 712
rect -35 -712 35 -280
<< xpolyres >>
rect -35 -280 35 280
<< locali >>
rect -165 808 -69 842
rect 69 808 165 842
rect -165 746 -131 808
rect 131 746 165 808
rect -165 -808 -131 -746
rect 131 -808 165 -746
rect -165 -842 -69 -808
rect 69 -842 165 -808
<< viali >>
rect -19 297 19 694
rect -19 -694 19 -297
<< metal1 >>
rect -25 694 25 706
rect -25 297 -19 694
rect 19 297 25 694
rect -25 285 25 297
rect -25 -297 25 -285
rect -25 -694 -19 -297
rect 19 -694 25 -297
rect -25 -706 25 -694
<< properties >>
string FIXED_BBOX -148 -825 148 825
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2.96 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 17.989k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
