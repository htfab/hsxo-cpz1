magic
tech sky130A
magscale 1 2
timestamp 1713747467
<< nwell >>
rect -2757 -3497 2757 3497
<< mvpmos >>
rect -2499 -3200 -2399 3200
rect -2341 -3200 -2241 3200
rect -2183 -3200 -2083 3200
rect -2025 -3200 -1925 3200
rect -1867 -3200 -1767 3200
rect -1709 -3200 -1609 3200
rect -1551 -3200 -1451 3200
rect -1393 -3200 -1293 3200
rect -1235 -3200 -1135 3200
rect -1077 -3200 -977 3200
rect -919 -3200 -819 3200
rect -761 -3200 -661 3200
rect -603 -3200 -503 3200
rect -445 -3200 -345 3200
rect -287 -3200 -187 3200
rect -129 -3200 -29 3200
rect 29 -3200 129 3200
rect 187 -3200 287 3200
rect 345 -3200 445 3200
rect 503 -3200 603 3200
rect 661 -3200 761 3200
rect 819 -3200 919 3200
rect 977 -3200 1077 3200
rect 1135 -3200 1235 3200
rect 1293 -3200 1393 3200
rect 1451 -3200 1551 3200
rect 1609 -3200 1709 3200
rect 1767 -3200 1867 3200
rect 1925 -3200 2025 3200
rect 2083 -3200 2183 3200
rect 2241 -3200 2341 3200
rect 2399 -3200 2499 3200
<< mvpdiff >>
rect -2557 3188 -2499 3200
rect -2557 -3188 -2545 3188
rect -2511 -3188 -2499 3188
rect -2557 -3200 -2499 -3188
rect -2399 3188 -2341 3200
rect -2399 -3188 -2387 3188
rect -2353 -3188 -2341 3188
rect -2399 -3200 -2341 -3188
rect -2241 3188 -2183 3200
rect -2241 -3188 -2229 3188
rect -2195 -3188 -2183 3188
rect -2241 -3200 -2183 -3188
rect -2083 3188 -2025 3200
rect -2083 -3188 -2071 3188
rect -2037 -3188 -2025 3188
rect -2083 -3200 -2025 -3188
rect -1925 3188 -1867 3200
rect -1925 -3188 -1913 3188
rect -1879 -3188 -1867 3188
rect -1925 -3200 -1867 -3188
rect -1767 3188 -1709 3200
rect -1767 -3188 -1755 3188
rect -1721 -3188 -1709 3188
rect -1767 -3200 -1709 -3188
rect -1609 3188 -1551 3200
rect -1609 -3188 -1597 3188
rect -1563 -3188 -1551 3188
rect -1609 -3200 -1551 -3188
rect -1451 3188 -1393 3200
rect -1451 -3188 -1439 3188
rect -1405 -3188 -1393 3188
rect -1451 -3200 -1393 -3188
rect -1293 3188 -1235 3200
rect -1293 -3188 -1281 3188
rect -1247 -3188 -1235 3188
rect -1293 -3200 -1235 -3188
rect -1135 3188 -1077 3200
rect -1135 -3188 -1123 3188
rect -1089 -3188 -1077 3188
rect -1135 -3200 -1077 -3188
rect -977 3188 -919 3200
rect -977 -3188 -965 3188
rect -931 -3188 -919 3188
rect -977 -3200 -919 -3188
rect -819 3188 -761 3200
rect -819 -3188 -807 3188
rect -773 -3188 -761 3188
rect -819 -3200 -761 -3188
rect -661 3188 -603 3200
rect -661 -3188 -649 3188
rect -615 -3188 -603 3188
rect -661 -3200 -603 -3188
rect -503 3188 -445 3200
rect -503 -3188 -491 3188
rect -457 -3188 -445 3188
rect -503 -3200 -445 -3188
rect -345 3188 -287 3200
rect -345 -3188 -333 3188
rect -299 -3188 -287 3188
rect -345 -3200 -287 -3188
rect -187 3188 -129 3200
rect -187 -3188 -175 3188
rect -141 -3188 -129 3188
rect -187 -3200 -129 -3188
rect -29 3188 29 3200
rect -29 -3188 -17 3188
rect 17 -3188 29 3188
rect -29 -3200 29 -3188
rect 129 3188 187 3200
rect 129 -3188 141 3188
rect 175 -3188 187 3188
rect 129 -3200 187 -3188
rect 287 3188 345 3200
rect 287 -3188 299 3188
rect 333 -3188 345 3188
rect 287 -3200 345 -3188
rect 445 3188 503 3200
rect 445 -3188 457 3188
rect 491 -3188 503 3188
rect 445 -3200 503 -3188
rect 603 3188 661 3200
rect 603 -3188 615 3188
rect 649 -3188 661 3188
rect 603 -3200 661 -3188
rect 761 3188 819 3200
rect 761 -3188 773 3188
rect 807 -3188 819 3188
rect 761 -3200 819 -3188
rect 919 3188 977 3200
rect 919 -3188 931 3188
rect 965 -3188 977 3188
rect 919 -3200 977 -3188
rect 1077 3188 1135 3200
rect 1077 -3188 1089 3188
rect 1123 -3188 1135 3188
rect 1077 -3200 1135 -3188
rect 1235 3188 1293 3200
rect 1235 -3188 1247 3188
rect 1281 -3188 1293 3188
rect 1235 -3200 1293 -3188
rect 1393 3188 1451 3200
rect 1393 -3188 1405 3188
rect 1439 -3188 1451 3188
rect 1393 -3200 1451 -3188
rect 1551 3188 1609 3200
rect 1551 -3188 1563 3188
rect 1597 -3188 1609 3188
rect 1551 -3200 1609 -3188
rect 1709 3188 1767 3200
rect 1709 -3188 1721 3188
rect 1755 -3188 1767 3188
rect 1709 -3200 1767 -3188
rect 1867 3188 1925 3200
rect 1867 -3188 1879 3188
rect 1913 -3188 1925 3188
rect 1867 -3200 1925 -3188
rect 2025 3188 2083 3200
rect 2025 -3188 2037 3188
rect 2071 -3188 2083 3188
rect 2025 -3200 2083 -3188
rect 2183 3188 2241 3200
rect 2183 -3188 2195 3188
rect 2229 -3188 2241 3188
rect 2183 -3200 2241 -3188
rect 2341 3188 2399 3200
rect 2341 -3188 2353 3188
rect 2387 -3188 2399 3188
rect 2341 -3200 2399 -3188
rect 2499 3188 2557 3200
rect 2499 -3188 2511 3188
rect 2545 -3188 2557 3188
rect 2499 -3200 2557 -3188
<< mvpdiffc >>
rect -2545 -3188 -2511 3188
rect -2387 -3188 -2353 3188
rect -2229 -3188 -2195 3188
rect -2071 -3188 -2037 3188
rect -1913 -3188 -1879 3188
rect -1755 -3188 -1721 3188
rect -1597 -3188 -1563 3188
rect -1439 -3188 -1405 3188
rect -1281 -3188 -1247 3188
rect -1123 -3188 -1089 3188
rect -965 -3188 -931 3188
rect -807 -3188 -773 3188
rect -649 -3188 -615 3188
rect -491 -3188 -457 3188
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
rect 457 -3188 491 3188
rect 615 -3188 649 3188
rect 773 -3188 807 3188
rect 931 -3188 965 3188
rect 1089 -3188 1123 3188
rect 1247 -3188 1281 3188
rect 1405 -3188 1439 3188
rect 1563 -3188 1597 3188
rect 1721 -3188 1755 3188
rect 1879 -3188 1913 3188
rect 2037 -3188 2071 3188
rect 2195 -3188 2229 3188
rect 2353 -3188 2387 3188
rect 2511 -3188 2545 3188
<< mvnsubdiff >>
rect -2691 3419 2691 3431
rect -2691 3385 -2583 3419
rect 2583 3385 2691 3419
rect -2691 3373 2691 3385
rect -2691 3323 -2633 3373
rect -2691 -3323 -2679 3323
rect -2645 -3323 -2633 3323
rect 2633 3323 2691 3373
rect -2691 -3373 -2633 -3323
rect 2633 -3323 2645 3323
rect 2679 -3323 2691 3323
rect 2633 -3373 2691 -3323
rect -2691 -3385 2691 -3373
rect -2691 -3419 -2583 -3385
rect 2583 -3419 2691 -3385
rect -2691 -3431 2691 -3419
<< mvnsubdiffcont >>
rect -2583 3385 2583 3419
rect -2679 -3323 -2645 3323
rect 2645 -3323 2679 3323
rect -2583 -3419 2583 -3385
<< poly >>
rect -2499 3281 -2399 3297
rect -2499 3247 -2483 3281
rect -2415 3247 -2399 3281
rect -2499 3200 -2399 3247
rect -2341 3281 -2241 3297
rect -2341 3247 -2325 3281
rect -2257 3247 -2241 3281
rect -2341 3200 -2241 3247
rect -2183 3281 -2083 3297
rect -2183 3247 -2167 3281
rect -2099 3247 -2083 3281
rect -2183 3200 -2083 3247
rect -2025 3281 -1925 3297
rect -2025 3247 -2009 3281
rect -1941 3247 -1925 3281
rect -2025 3200 -1925 3247
rect -1867 3281 -1767 3297
rect -1867 3247 -1851 3281
rect -1783 3247 -1767 3281
rect -1867 3200 -1767 3247
rect -1709 3281 -1609 3297
rect -1709 3247 -1693 3281
rect -1625 3247 -1609 3281
rect -1709 3200 -1609 3247
rect -1551 3281 -1451 3297
rect -1551 3247 -1535 3281
rect -1467 3247 -1451 3281
rect -1551 3200 -1451 3247
rect -1393 3281 -1293 3297
rect -1393 3247 -1377 3281
rect -1309 3247 -1293 3281
rect -1393 3200 -1293 3247
rect -1235 3281 -1135 3297
rect -1235 3247 -1219 3281
rect -1151 3247 -1135 3281
rect -1235 3200 -1135 3247
rect -1077 3281 -977 3297
rect -1077 3247 -1061 3281
rect -993 3247 -977 3281
rect -1077 3200 -977 3247
rect -919 3281 -819 3297
rect -919 3247 -903 3281
rect -835 3247 -819 3281
rect -919 3200 -819 3247
rect -761 3281 -661 3297
rect -761 3247 -745 3281
rect -677 3247 -661 3281
rect -761 3200 -661 3247
rect -603 3281 -503 3297
rect -603 3247 -587 3281
rect -519 3247 -503 3281
rect -603 3200 -503 3247
rect -445 3281 -345 3297
rect -445 3247 -429 3281
rect -361 3247 -345 3281
rect -445 3200 -345 3247
rect -287 3281 -187 3297
rect -287 3247 -271 3281
rect -203 3247 -187 3281
rect -287 3200 -187 3247
rect -129 3281 -29 3297
rect -129 3247 -113 3281
rect -45 3247 -29 3281
rect -129 3200 -29 3247
rect 29 3281 129 3297
rect 29 3247 45 3281
rect 113 3247 129 3281
rect 29 3200 129 3247
rect 187 3281 287 3297
rect 187 3247 203 3281
rect 271 3247 287 3281
rect 187 3200 287 3247
rect 345 3281 445 3297
rect 345 3247 361 3281
rect 429 3247 445 3281
rect 345 3200 445 3247
rect 503 3281 603 3297
rect 503 3247 519 3281
rect 587 3247 603 3281
rect 503 3200 603 3247
rect 661 3281 761 3297
rect 661 3247 677 3281
rect 745 3247 761 3281
rect 661 3200 761 3247
rect 819 3281 919 3297
rect 819 3247 835 3281
rect 903 3247 919 3281
rect 819 3200 919 3247
rect 977 3281 1077 3297
rect 977 3247 993 3281
rect 1061 3247 1077 3281
rect 977 3200 1077 3247
rect 1135 3281 1235 3297
rect 1135 3247 1151 3281
rect 1219 3247 1235 3281
rect 1135 3200 1235 3247
rect 1293 3281 1393 3297
rect 1293 3247 1309 3281
rect 1377 3247 1393 3281
rect 1293 3200 1393 3247
rect 1451 3281 1551 3297
rect 1451 3247 1467 3281
rect 1535 3247 1551 3281
rect 1451 3200 1551 3247
rect 1609 3281 1709 3297
rect 1609 3247 1625 3281
rect 1693 3247 1709 3281
rect 1609 3200 1709 3247
rect 1767 3281 1867 3297
rect 1767 3247 1783 3281
rect 1851 3247 1867 3281
rect 1767 3200 1867 3247
rect 1925 3281 2025 3297
rect 1925 3247 1941 3281
rect 2009 3247 2025 3281
rect 1925 3200 2025 3247
rect 2083 3281 2183 3297
rect 2083 3247 2099 3281
rect 2167 3247 2183 3281
rect 2083 3200 2183 3247
rect 2241 3281 2341 3297
rect 2241 3247 2257 3281
rect 2325 3247 2341 3281
rect 2241 3200 2341 3247
rect 2399 3281 2499 3297
rect 2399 3247 2415 3281
rect 2483 3247 2499 3281
rect 2399 3200 2499 3247
rect -2499 -3247 -2399 -3200
rect -2499 -3281 -2483 -3247
rect -2415 -3281 -2399 -3247
rect -2499 -3297 -2399 -3281
rect -2341 -3247 -2241 -3200
rect -2341 -3281 -2325 -3247
rect -2257 -3281 -2241 -3247
rect -2341 -3297 -2241 -3281
rect -2183 -3247 -2083 -3200
rect -2183 -3281 -2167 -3247
rect -2099 -3281 -2083 -3247
rect -2183 -3297 -2083 -3281
rect -2025 -3247 -1925 -3200
rect -2025 -3281 -2009 -3247
rect -1941 -3281 -1925 -3247
rect -2025 -3297 -1925 -3281
rect -1867 -3247 -1767 -3200
rect -1867 -3281 -1851 -3247
rect -1783 -3281 -1767 -3247
rect -1867 -3297 -1767 -3281
rect -1709 -3247 -1609 -3200
rect -1709 -3281 -1693 -3247
rect -1625 -3281 -1609 -3247
rect -1709 -3297 -1609 -3281
rect -1551 -3247 -1451 -3200
rect -1551 -3281 -1535 -3247
rect -1467 -3281 -1451 -3247
rect -1551 -3297 -1451 -3281
rect -1393 -3247 -1293 -3200
rect -1393 -3281 -1377 -3247
rect -1309 -3281 -1293 -3247
rect -1393 -3297 -1293 -3281
rect -1235 -3247 -1135 -3200
rect -1235 -3281 -1219 -3247
rect -1151 -3281 -1135 -3247
rect -1235 -3297 -1135 -3281
rect -1077 -3247 -977 -3200
rect -1077 -3281 -1061 -3247
rect -993 -3281 -977 -3247
rect -1077 -3297 -977 -3281
rect -919 -3247 -819 -3200
rect -919 -3281 -903 -3247
rect -835 -3281 -819 -3247
rect -919 -3297 -819 -3281
rect -761 -3247 -661 -3200
rect -761 -3281 -745 -3247
rect -677 -3281 -661 -3247
rect -761 -3297 -661 -3281
rect -603 -3247 -503 -3200
rect -603 -3281 -587 -3247
rect -519 -3281 -503 -3247
rect -603 -3297 -503 -3281
rect -445 -3247 -345 -3200
rect -445 -3281 -429 -3247
rect -361 -3281 -345 -3247
rect -445 -3297 -345 -3281
rect -287 -3247 -187 -3200
rect -287 -3281 -271 -3247
rect -203 -3281 -187 -3247
rect -287 -3297 -187 -3281
rect -129 -3247 -29 -3200
rect -129 -3281 -113 -3247
rect -45 -3281 -29 -3247
rect -129 -3297 -29 -3281
rect 29 -3247 129 -3200
rect 29 -3281 45 -3247
rect 113 -3281 129 -3247
rect 29 -3297 129 -3281
rect 187 -3247 287 -3200
rect 187 -3281 203 -3247
rect 271 -3281 287 -3247
rect 187 -3297 287 -3281
rect 345 -3247 445 -3200
rect 345 -3281 361 -3247
rect 429 -3281 445 -3247
rect 345 -3297 445 -3281
rect 503 -3247 603 -3200
rect 503 -3281 519 -3247
rect 587 -3281 603 -3247
rect 503 -3297 603 -3281
rect 661 -3247 761 -3200
rect 661 -3281 677 -3247
rect 745 -3281 761 -3247
rect 661 -3297 761 -3281
rect 819 -3247 919 -3200
rect 819 -3281 835 -3247
rect 903 -3281 919 -3247
rect 819 -3297 919 -3281
rect 977 -3247 1077 -3200
rect 977 -3281 993 -3247
rect 1061 -3281 1077 -3247
rect 977 -3297 1077 -3281
rect 1135 -3247 1235 -3200
rect 1135 -3281 1151 -3247
rect 1219 -3281 1235 -3247
rect 1135 -3297 1235 -3281
rect 1293 -3247 1393 -3200
rect 1293 -3281 1309 -3247
rect 1377 -3281 1393 -3247
rect 1293 -3297 1393 -3281
rect 1451 -3247 1551 -3200
rect 1451 -3281 1467 -3247
rect 1535 -3281 1551 -3247
rect 1451 -3297 1551 -3281
rect 1609 -3247 1709 -3200
rect 1609 -3281 1625 -3247
rect 1693 -3281 1709 -3247
rect 1609 -3297 1709 -3281
rect 1767 -3247 1867 -3200
rect 1767 -3281 1783 -3247
rect 1851 -3281 1867 -3247
rect 1767 -3297 1867 -3281
rect 1925 -3247 2025 -3200
rect 1925 -3281 1941 -3247
rect 2009 -3281 2025 -3247
rect 1925 -3297 2025 -3281
rect 2083 -3247 2183 -3200
rect 2083 -3281 2099 -3247
rect 2167 -3281 2183 -3247
rect 2083 -3297 2183 -3281
rect 2241 -3247 2341 -3200
rect 2241 -3281 2257 -3247
rect 2325 -3281 2341 -3247
rect 2241 -3297 2341 -3281
rect 2399 -3247 2499 -3200
rect 2399 -3281 2415 -3247
rect 2483 -3281 2499 -3247
rect 2399 -3297 2499 -3281
<< polycont >>
rect -2483 3247 -2415 3281
rect -2325 3247 -2257 3281
rect -2167 3247 -2099 3281
rect -2009 3247 -1941 3281
rect -1851 3247 -1783 3281
rect -1693 3247 -1625 3281
rect -1535 3247 -1467 3281
rect -1377 3247 -1309 3281
rect -1219 3247 -1151 3281
rect -1061 3247 -993 3281
rect -903 3247 -835 3281
rect -745 3247 -677 3281
rect -587 3247 -519 3281
rect -429 3247 -361 3281
rect -271 3247 -203 3281
rect -113 3247 -45 3281
rect 45 3247 113 3281
rect 203 3247 271 3281
rect 361 3247 429 3281
rect 519 3247 587 3281
rect 677 3247 745 3281
rect 835 3247 903 3281
rect 993 3247 1061 3281
rect 1151 3247 1219 3281
rect 1309 3247 1377 3281
rect 1467 3247 1535 3281
rect 1625 3247 1693 3281
rect 1783 3247 1851 3281
rect 1941 3247 2009 3281
rect 2099 3247 2167 3281
rect 2257 3247 2325 3281
rect 2415 3247 2483 3281
rect -2483 -3281 -2415 -3247
rect -2325 -3281 -2257 -3247
rect -2167 -3281 -2099 -3247
rect -2009 -3281 -1941 -3247
rect -1851 -3281 -1783 -3247
rect -1693 -3281 -1625 -3247
rect -1535 -3281 -1467 -3247
rect -1377 -3281 -1309 -3247
rect -1219 -3281 -1151 -3247
rect -1061 -3281 -993 -3247
rect -903 -3281 -835 -3247
rect -745 -3281 -677 -3247
rect -587 -3281 -519 -3247
rect -429 -3281 -361 -3247
rect -271 -3281 -203 -3247
rect -113 -3281 -45 -3247
rect 45 -3281 113 -3247
rect 203 -3281 271 -3247
rect 361 -3281 429 -3247
rect 519 -3281 587 -3247
rect 677 -3281 745 -3247
rect 835 -3281 903 -3247
rect 993 -3281 1061 -3247
rect 1151 -3281 1219 -3247
rect 1309 -3281 1377 -3247
rect 1467 -3281 1535 -3247
rect 1625 -3281 1693 -3247
rect 1783 -3281 1851 -3247
rect 1941 -3281 2009 -3247
rect 2099 -3281 2167 -3247
rect 2257 -3281 2325 -3247
rect 2415 -3281 2483 -3247
<< locali >>
rect -2679 3385 -2583 3419
rect 2583 3385 2679 3419
rect -2679 3323 -2645 3385
rect 2645 3323 2679 3385
rect -2499 3247 -2483 3281
rect -2415 3247 -2399 3281
rect -2341 3247 -2325 3281
rect -2257 3247 -2241 3281
rect -2183 3247 -2167 3281
rect -2099 3247 -2083 3281
rect -2025 3247 -2009 3281
rect -1941 3247 -1925 3281
rect -1867 3247 -1851 3281
rect -1783 3247 -1767 3281
rect -1709 3247 -1693 3281
rect -1625 3247 -1609 3281
rect -1551 3247 -1535 3281
rect -1467 3247 -1451 3281
rect -1393 3247 -1377 3281
rect -1309 3247 -1293 3281
rect -1235 3247 -1219 3281
rect -1151 3247 -1135 3281
rect -1077 3247 -1061 3281
rect -993 3247 -977 3281
rect -919 3247 -903 3281
rect -835 3247 -819 3281
rect -761 3247 -745 3281
rect -677 3247 -661 3281
rect -603 3247 -587 3281
rect -519 3247 -503 3281
rect -445 3247 -429 3281
rect -361 3247 -345 3281
rect -287 3247 -271 3281
rect -203 3247 -187 3281
rect -129 3247 -113 3281
rect -45 3247 -29 3281
rect 29 3247 45 3281
rect 113 3247 129 3281
rect 187 3247 203 3281
rect 271 3247 287 3281
rect 345 3247 361 3281
rect 429 3247 445 3281
rect 503 3247 519 3281
rect 587 3247 603 3281
rect 661 3247 677 3281
rect 745 3247 761 3281
rect 819 3247 835 3281
rect 903 3247 919 3281
rect 977 3247 993 3281
rect 1061 3247 1077 3281
rect 1135 3247 1151 3281
rect 1219 3247 1235 3281
rect 1293 3247 1309 3281
rect 1377 3247 1393 3281
rect 1451 3247 1467 3281
rect 1535 3247 1551 3281
rect 1609 3247 1625 3281
rect 1693 3247 1709 3281
rect 1767 3247 1783 3281
rect 1851 3247 1867 3281
rect 1925 3247 1941 3281
rect 2009 3247 2025 3281
rect 2083 3247 2099 3281
rect 2167 3247 2183 3281
rect 2241 3247 2257 3281
rect 2325 3247 2341 3281
rect 2399 3247 2415 3281
rect 2483 3247 2499 3281
rect -2545 3188 -2511 3204
rect -2545 -3204 -2511 -3188
rect -2387 3188 -2353 3204
rect -2387 -3204 -2353 -3188
rect -2229 3188 -2195 3204
rect -2229 -3204 -2195 -3188
rect -2071 3188 -2037 3204
rect -2071 -3204 -2037 -3188
rect -1913 3188 -1879 3204
rect -1913 -3204 -1879 -3188
rect -1755 3188 -1721 3204
rect -1755 -3204 -1721 -3188
rect -1597 3188 -1563 3204
rect -1597 -3204 -1563 -3188
rect -1439 3188 -1405 3204
rect -1439 -3204 -1405 -3188
rect -1281 3188 -1247 3204
rect -1281 -3204 -1247 -3188
rect -1123 3188 -1089 3204
rect -1123 -3204 -1089 -3188
rect -965 3188 -931 3204
rect -965 -3204 -931 -3188
rect -807 3188 -773 3204
rect -807 -3204 -773 -3188
rect -649 3188 -615 3204
rect -649 -3204 -615 -3188
rect -491 3188 -457 3204
rect -491 -3204 -457 -3188
rect -333 3188 -299 3204
rect -333 -3204 -299 -3188
rect -175 3188 -141 3204
rect -175 -3204 -141 -3188
rect -17 3188 17 3204
rect -17 -3204 17 -3188
rect 141 3188 175 3204
rect 141 -3204 175 -3188
rect 299 3188 333 3204
rect 299 -3204 333 -3188
rect 457 3188 491 3204
rect 457 -3204 491 -3188
rect 615 3188 649 3204
rect 615 -3204 649 -3188
rect 773 3188 807 3204
rect 773 -3204 807 -3188
rect 931 3188 965 3204
rect 931 -3204 965 -3188
rect 1089 3188 1123 3204
rect 1089 -3204 1123 -3188
rect 1247 3188 1281 3204
rect 1247 -3204 1281 -3188
rect 1405 3188 1439 3204
rect 1405 -3204 1439 -3188
rect 1563 3188 1597 3204
rect 1563 -3204 1597 -3188
rect 1721 3188 1755 3204
rect 1721 -3204 1755 -3188
rect 1879 3188 1913 3204
rect 1879 -3204 1913 -3188
rect 2037 3188 2071 3204
rect 2037 -3204 2071 -3188
rect 2195 3188 2229 3204
rect 2195 -3204 2229 -3188
rect 2353 3188 2387 3204
rect 2353 -3204 2387 -3188
rect 2511 3188 2545 3204
rect 2511 -3204 2545 -3188
rect -2499 -3281 -2483 -3247
rect -2415 -3281 -2399 -3247
rect -2341 -3281 -2325 -3247
rect -2257 -3281 -2241 -3247
rect -2183 -3281 -2167 -3247
rect -2099 -3281 -2083 -3247
rect -2025 -3281 -2009 -3247
rect -1941 -3281 -1925 -3247
rect -1867 -3281 -1851 -3247
rect -1783 -3281 -1767 -3247
rect -1709 -3281 -1693 -3247
rect -1625 -3281 -1609 -3247
rect -1551 -3281 -1535 -3247
rect -1467 -3281 -1451 -3247
rect -1393 -3281 -1377 -3247
rect -1309 -3281 -1293 -3247
rect -1235 -3281 -1219 -3247
rect -1151 -3281 -1135 -3247
rect -1077 -3281 -1061 -3247
rect -993 -3281 -977 -3247
rect -919 -3281 -903 -3247
rect -835 -3281 -819 -3247
rect -761 -3281 -745 -3247
rect -677 -3281 -661 -3247
rect -603 -3281 -587 -3247
rect -519 -3281 -503 -3247
rect -445 -3281 -429 -3247
rect -361 -3281 -345 -3247
rect -287 -3281 -271 -3247
rect -203 -3281 -187 -3247
rect -129 -3281 -113 -3247
rect -45 -3281 -29 -3247
rect 29 -3281 45 -3247
rect 113 -3281 129 -3247
rect 187 -3281 203 -3247
rect 271 -3281 287 -3247
rect 345 -3281 361 -3247
rect 429 -3281 445 -3247
rect 503 -3281 519 -3247
rect 587 -3281 603 -3247
rect 661 -3281 677 -3247
rect 745 -3281 761 -3247
rect 819 -3281 835 -3247
rect 903 -3281 919 -3247
rect 977 -3281 993 -3247
rect 1061 -3281 1077 -3247
rect 1135 -3281 1151 -3247
rect 1219 -3281 1235 -3247
rect 1293 -3281 1309 -3247
rect 1377 -3281 1393 -3247
rect 1451 -3281 1467 -3247
rect 1535 -3281 1551 -3247
rect 1609 -3281 1625 -3247
rect 1693 -3281 1709 -3247
rect 1767 -3281 1783 -3247
rect 1851 -3281 1867 -3247
rect 1925 -3281 1941 -3247
rect 2009 -3281 2025 -3247
rect 2083 -3281 2099 -3247
rect 2167 -3281 2183 -3247
rect 2241 -3281 2257 -3247
rect 2325 -3281 2341 -3247
rect 2399 -3281 2415 -3247
rect 2483 -3281 2499 -3247
rect -2679 -3385 -2645 -3323
rect 2645 -3385 2679 -3323
rect -2679 -3419 -2583 -3385
rect 2583 -3419 2679 -3385
<< viali >>
rect -2483 3247 -2415 3281
rect -2325 3247 -2257 3281
rect -2167 3247 -2099 3281
rect -2009 3247 -1941 3281
rect -1851 3247 -1783 3281
rect -1693 3247 -1625 3281
rect -1535 3247 -1467 3281
rect -1377 3247 -1309 3281
rect -1219 3247 -1151 3281
rect -1061 3247 -993 3281
rect -903 3247 -835 3281
rect -745 3247 -677 3281
rect -587 3247 -519 3281
rect -429 3247 -361 3281
rect -271 3247 -203 3281
rect -113 3247 -45 3281
rect 45 3247 113 3281
rect 203 3247 271 3281
rect 361 3247 429 3281
rect 519 3247 587 3281
rect 677 3247 745 3281
rect 835 3247 903 3281
rect 993 3247 1061 3281
rect 1151 3247 1219 3281
rect 1309 3247 1377 3281
rect 1467 3247 1535 3281
rect 1625 3247 1693 3281
rect 1783 3247 1851 3281
rect 1941 3247 2009 3281
rect 2099 3247 2167 3281
rect 2257 3247 2325 3281
rect 2415 3247 2483 3281
rect -2545 -3188 -2511 3188
rect -2387 -3188 -2353 3188
rect -2229 -3188 -2195 3188
rect -2071 -3188 -2037 3188
rect -1913 -3188 -1879 3188
rect -1755 -3188 -1721 3188
rect -1597 -3188 -1563 3188
rect -1439 -3188 -1405 3188
rect -1281 -3188 -1247 3188
rect -1123 -3188 -1089 3188
rect -965 -3188 -931 3188
rect -807 -3188 -773 3188
rect -649 -3188 -615 3188
rect -491 -3188 -457 3188
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
rect 457 -3188 491 3188
rect 615 -3188 649 3188
rect 773 -3188 807 3188
rect 931 -3188 965 3188
rect 1089 -3188 1123 3188
rect 1247 -3188 1281 3188
rect 1405 -3188 1439 3188
rect 1563 -3188 1597 3188
rect 1721 -3188 1755 3188
rect 1879 -3188 1913 3188
rect 2037 -3188 2071 3188
rect 2195 -3188 2229 3188
rect 2353 -3188 2387 3188
rect 2511 -3188 2545 3188
rect -2483 -3281 -2415 -3247
rect -2325 -3281 -2257 -3247
rect -2167 -3281 -2099 -3247
rect -2009 -3281 -1941 -3247
rect -1851 -3281 -1783 -3247
rect -1693 -3281 -1625 -3247
rect -1535 -3281 -1467 -3247
rect -1377 -3281 -1309 -3247
rect -1219 -3281 -1151 -3247
rect -1061 -3281 -993 -3247
rect -903 -3281 -835 -3247
rect -745 -3281 -677 -3247
rect -587 -3281 -519 -3247
rect -429 -3281 -361 -3247
rect -271 -3281 -203 -3247
rect -113 -3281 -45 -3247
rect 45 -3281 113 -3247
rect 203 -3281 271 -3247
rect 361 -3281 429 -3247
rect 519 -3281 587 -3247
rect 677 -3281 745 -3247
rect 835 -3281 903 -3247
rect 993 -3281 1061 -3247
rect 1151 -3281 1219 -3247
rect 1309 -3281 1377 -3247
rect 1467 -3281 1535 -3247
rect 1625 -3281 1693 -3247
rect 1783 -3281 1851 -3247
rect 1941 -3281 2009 -3247
rect 2099 -3281 2167 -3247
rect 2257 -3281 2325 -3247
rect 2415 -3281 2483 -3247
<< metal1 >>
rect -2495 3281 -2403 3287
rect -2495 3247 -2483 3281
rect -2415 3247 -2403 3281
rect -2495 3241 -2403 3247
rect -2337 3281 -2245 3287
rect -2337 3247 -2325 3281
rect -2257 3247 -2245 3281
rect -2337 3241 -2245 3247
rect -2179 3281 -2087 3287
rect -2179 3247 -2167 3281
rect -2099 3247 -2087 3281
rect -2179 3241 -2087 3247
rect -2021 3281 -1929 3287
rect -2021 3247 -2009 3281
rect -1941 3247 -1929 3281
rect -2021 3241 -1929 3247
rect -1863 3281 -1771 3287
rect -1863 3247 -1851 3281
rect -1783 3247 -1771 3281
rect -1863 3241 -1771 3247
rect -1705 3281 -1613 3287
rect -1705 3247 -1693 3281
rect -1625 3247 -1613 3281
rect -1705 3241 -1613 3247
rect -1547 3281 -1455 3287
rect -1547 3247 -1535 3281
rect -1467 3247 -1455 3281
rect -1547 3241 -1455 3247
rect -1389 3281 -1297 3287
rect -1389 3247 -1377 3281
rect -1309 3247 -1297 3281
rect -1389 3241 -1297 3247
rect -1231 3281 -1139 3287
rect -1231 3247 -1219 3281
rect -1151 3247 -1139 3281
rect -1231 3241 -1139 3247
rect -1073 3281 -981 3287
rect -1073 3247 -1061 3281
rect -993 3247 -981 3281
rect -1073 3241 -981 3247
rect -915 3281 -823 3287
rect -915 3247 -903 3281
rect -835 3247 -823 3281
rect -915 3241 -823 3247
rect -757 3281 -665 3287
rect -757 3247 -745 3281
rect -677 3247 -665 3281
rect -757 3241 -665 3247
rect -599 3281 -507 3287
rect -599 3247 -587 3281
rect -519 3247 -507 3281
rect -599 3241 -507 3247
rect -441 3281 -349 3287
rect -441 3247 -429 3281
rect -361 3247 -349 3281
rect -441 3241 -349 3247
rect -283 3281 -191 3287
rect -283 3247 -271 3281
rect -203 3247 -191 3281
rect -283 3241 -191 3247
rect -125 3281 -33 3287
rect -125 3247 -113 3281
rect -45 3247 -33 3281
rect -125 3241 -33 3247
rect 33 3281 125 3287
rect 33 3247 45 3281
rect 113 3247 125 3281
rect 33 3241 125 3247
rect 191 3281 283 3287
rect 191 3247 203 3281
rect 271 3247 283 3281
rect 191 3241 283 3247
rect 349 3281 441 3287
rect 349 3247 361 3281
rect 429 3247 441 3281
rect 349 3241 441 3247
rect 507 3281 599 3287
rect 507 3247 519 3281
rect 587 3247 599 3281
rect 507 3241 599 3247
rect 665 3281 757 3287
rect 665 3247 677 3281
rect 745 3247 757 3281
rect 665 3241 757 3247
rect 823 3281 915 3287
rect 823 3247 835 3281
rect 903 3247 915 3281
rect 823 3241 915 3247
rect 981 3281 1073 3287
rect 981 3247 993 3281
rect 1061 3247 1073 3281
rect 981 3241 1073 3247
rect 1139 3281 1231 3287
rect 1139 3247 1151 3281
rect 1219 3247 1231 3281
rect 1139 3241 1231 3247
rect 1297 3281 1389 3287
rect 1297 3247 1309 3281
rect 1377 3247 1389 3281
rect 1297 3241 1389 3247
rect 1455 3281 1547 3287
rect 1455 3247 1467 3281
rect 1535 3247 1547 3281
rect 1455 3241 1547 3247
rect 1613 3281 1705 3287
rect 1613 3247 1625 3281
rect 1693 3247 1705 3281
rect 1613 3241 1705 3247
rect 1771 3281 1863 3287
rect 1771 3247 1783 3281
rect 1851 3247 1863 3281
rect 1771 3241 1863 3247
rect 1929 3281 2021 3287
rect 1929 3247 1941 3281
rect 2009 3247 2021 3281
rect 1929 3241 2021 3247
rect 2087 3281 2179 3287
rect 2087 3247 2099 3281
rect 2167 3247 2179 3281
rect 2087 3241 2179 3247
rect 2245 3281 2337 3287
rect 2245 3247 2257 3281
rect 2325 3247 2337 3281
rect 2245 3241 2337 3247
rect 2403 3281 2495 3287
rect 2403 3247 2415 3281
rect 2483 3247 2495 3281
rect 2403 3241 2495 3247
rect -2551 3188 -2505 3200
rect -2551 -3188 -2545 3188
rect -2511 -3188 -2505 3188
rect -2551 -3200 -2505 -3188
rect -2393 3188 -2347 3200
rect -2393 -3188 -2387 3188
rect -2353 -3188 -2347 3188
rect -2393 -3200 -2347 -3188
rect -2235 3188 -2189 3200
rect -2235 -3188 -2229 3188
rect -2195 -3188 -2189 3188
rect -2235 -3200 -2189 -3188
rect -2077 3188 -2031 3200
rect -2077 -3188 -2071 3188
rect -2037 -3188 -2031 3188
rect -2077 -3200 -2031 -3188
rect -1919 3188 -1873 3200
rect -1919 -3188 -1913 3188
rect -1879 -3188 -1873 3188
rect -1919 -3200 -1873 -3188
rect -1761 3188 -1715 3200
rect -1761 -3188 -1755 3188
rect -1721 -3188 -1715 3188
rect -1761 -3200 -1715 -3188
rect -1603 3188 -1557 3200
rect -1603 -3188 -1597 3188
rect -1563 -3188 -1557 3188
rect -1603 -3200 -1557 -3188
rect -1445 3188 -1399 3200
rect -1445 -3188 -1439 3188
rect -1405 -3188 -1399 3188
rect -1445 -3200 -1399 -3188
rect -1287 3188 -1241 3200
rect -1287 -3188 -1281 3188
rect -1247 -3188 -1241 3188
rect -1287 -3200 -1241 -3188
rect -1129 3188 -1083 3200
rect -1129 -3188 -1123 3188
rect -1089 -3188 -1083 3188
rect -1129 -3200 -1083 -3188
rect -971 3188 -925 3200
rect -971 -3188 -965 3188
rect -931 -3188 -925 3188
rect -971 -3200 -925 -3188
rect -813 3188 -767 3200
rect -813 -3188 -807 3188
rect -773 -3188 -767 3188
rect -813 -3200 -767 -3188
rect -655 3188 -609 3200
rect -655 -3188 -649 3188
rect -615 -3188 -609 3188
rect -655 -3200 -609 -3188
rect -497 3188 -451 3200
rect -497 -3188 -491 3188
rect -457 -3188 -451 3188
rect -497 -3200 -451 -3188
rect -339 3188 -293 3200
rect -339 -3188 -333 3188
rect -299 -3188 -293 3188
rect -339 -3200 -293 -3188
rect -181 3188 -135 3200
rect -181 -3188 -175 3188
rect -141 -3188 -135 3188
rect -181 -3200 -135 -3188
rect -23 3188 23 3200
rect -23 -3188 -17 3188
rect 17 -3188 23 3188
rect -23 -3200 23 -3188
rect 135 3188 181 3200
rect 135 -3188 141 3188
rect 175 -3188 181 3188
rect 135 -3200 181 -3188
rect 293 3188 339 3200
rect 293 -3188 299 3188
rect 333 -3188 339 3188
rect 293 -3200 339 -3188
rect 451 3188 497 3200
rect 451 -3188 457 3188
rect 491 -3188 497 3188
rect 451 -3200 497 -3188
rect 609 3188 655 3200
rect 609 -3188 615 3188
rect 649 -3188 655 3188
rect 609 -3200 655 -3188
rect 767 3188 813 3200
rect 767 -3188 773 3188
rect 807 -3188 813 3188
rect 767 -3200 813 -3188
rect 925 3188 971 3200
rect 925 -3188 931 3188
rect 965 -3188 971 3188
rect 925 -3200 971 -3188
rect 1083 3188 1129 3200
rect 1083 -3188 1089 3188
rect 1123 -3188 1129 3188
rect 1083 -3200 1129 -3188
rect 1241 3188 1287 3200
rect 1241 -3188 1247 3188
rect 1281 -3188 1287 3188
rect 1241 -3200 1287 -3188
rect 1399 3188 1445 3200
rect 1399 -3188 1405 3188
rect 1439 -3188 1445 3188
rect 1399 -3200 1445 -3188
rect 1557 3188 1603 3200
rect 1557 -3188 1563 3188
rect 1597 -3188 1603 3188
rect 1557 -3200 1603 -3188
rect 1715 3188 1761 3200
rect 1715 -3188 1721 3188
rect 1755 -3188 1761 3188
rect 1715 -3200 1761 -3188
rect 1873 3188 1919 3200
rect 1873 -3188 1879 3188
rect 1913 -3188 1919 3188
rect 1873 -3200 1919 -3188
rect 2031 3188 2077 3200
rect 2031 -3188 2037 3188
rect 2071 -3188 2077 3188
rect 2031 -3200 2077 -3188
rect 2189 3188 2235 3200
rect 2189 -3188 2195 3188
rect 2229 -3188 2235 3188
rect 2189 -3200 2235 -3188
rect 2347 3188 2393 3200
rect 2347 -3188 2353 3188
rect 2387 -3188 2393 3188
rect 2347 -3200 2393 -3188
rect 2505 3188 2551 3200
rect 2505 -3188 2511 3188
rect 2545 -3188 2551 3188
rect 2505 -3200 2551 -3188
rect -2495 -3247 -2403 -3241
rect -2495 -3281 -2483 -3247
rect -2415 -3281 -2403 -3247
rect -2495 -3287 -2403 -3281
rect -2337 -3247 -2245 -3241
rect -2337 -3281 -2325 -3247
rect -2257 -3281 -2245 -3247
rect -2337 -3287 -2245 -3281
rect -2179 -3247 -2087 -3241
rect -2179 -3281 -2167 -3247
rect -2099 -3281 -2087 -3247
rect -2179 -3287 -2087 -3281
rect -2021 -3247 -1929 -3241
rect -2021 -3281 -2009 -3247
rect -1941 -3281 -1929 -3247
rect -2021 -3287 -1929 -3281
rect -1863 -3247 -1771 -3241
rect -1863 -3281 -1851 -3247
rect -1783 -3281 -1771 -3247
rect -1863 -3287 -1771 -3281
rect -1705 -3247 -1613 -3241
rect -1705 -3281 -1693 -3247
rect -1625 -3281 -1613 -3247
rect -1705 -3287 -1613 -3281
rect -1547 -3247 -1455 -3241
rect -1547 -3281 -1535 -3247
rect -1467 -3281 -1455 -3247
rect -1547 -3287 -1455 -3281
rect -1389 -3247 -1297 -3241
rect -1389 -3281 -1377 -3247
rect -1309 -3281 -1297 -3247
rect -1389 -3287 -1297 -3281
rect -1231 -3247 -1139 -3241
rect -1231 -3281 -1219 -3247
rect -1151 -3281 -1139 -3247
rect -1231 -3287 -1139 -3281
rect -1073 -3247 -981 -3241
rect -1073 -3281 -1061 -3247
rect -993 -3281 -981 -3247
rect -1073 -3287 -981 -3281
rect -915 -3247 -823 -3241
rect -915 -3281 -903 -3247
rect -835 -3281 -823 -3247
rect -915 -3287 -823 -3281
rect -757 -3247 -665 -3241
rect -757 -3281 -745 -3247
rect -677 -3281 -665 -3247
rect -757 -3287 -665 -3281
rect -599 -3247 -507 -3241
rect -599 -3281 -587 -3247
rect -519 -3281 -507 -3247
rect -599 -3287 -507 -3281
rect -441 -3247 -349 -3241
rect -441 -3281 -429 -3247
rect -361 -3281 -349 -3247
rect -441 -3287 -349 -3281
rect -283 -3247 -191 -3241
rect -283 -3281 -271 -3247
rect -203 -3281 -191 -3247
rect -283 -3287 -191 -3281
rect -125 -3247 -33 -3241
rect -125 -3281 -113 -3247
rect -45 -3281 -33 -3247
rect -125 -3287 -33 -3281
rect 33 -3247 125 -3241
rect 33 -3281 45 -3247
rect 113 -3281 125 -3247
rect 33 -3287 125 -3281
rect 191 -3247 283 -3241
rect 191 -3281 203 -3247
rect 271 -3281 283 -3247
rect 191 -3287 283 -3281
rect 349 -3247 441 -3241
rect 349 -3281 361 -3247
rect 429 -3281 441 -3247
rect 349 -3287 441 -3281
rect 507 -3247 599 -3241
rect 507 -3281 519 -3247
rect 587 -3281 599 -3247
rect 507 -3287 599 -3281
rect 665 -3247 757 -3241
rect 665 -3281 677 -3247
rect 745 -3281 757 -3247
rect 665 -3287 757 -3281
rect 823 -3247 915 -3241
rect 823 -3281 835 -3247
rect 903 -3281 915 -3247
rect 823 -3287 915 -3281
rect 981 -3247 1073 -3241
rect 981 -3281 993 -3247
rect 1061 -3281 1073 -3247
rect 981 -3287 1073 -3281
rect 1139 -3247 1231 -3241
rect 1139 -3281 1151 -3247
rect 1219 -3281 1231 -3247
rect 1139 -3287 1231 -3281
rect 1297 -3247 1389 -3241
rect 1297 -3281 1309 -3247
rect 1377 -3281 1389 -3247
rect 1297 -3287 1389 -3281
rect 1455 -3247 1547 -3241
rect 1455 -3281 1467 -3247
rect 1535 -3281 1547 -3247
rect 1455 -3287 1547 -3281
rect 1613 -3247 1705 -3241
rect 1613 -3281 1625 -3247
rect 1693 -3281 1705 -3247
rect 1613 -3287 1705 -3281
rect 1771 -3247 1863 -3241
rect 1771 -3281 1783 -3247
rect 1851 -3281 1863 -3247
rect 1771 -3287 1863 -3281
rect 1929 -3247 2021 -3241
rect 1929 -3281 1941 -3247
rect 2009 -3281 2021 -3247
rect 1929 -3287 2021 -3281
rect 2087 -3247 2179 -3241
rect 2087 -3281 2099 -3247
rect 2167 -3281 2179 -3247
rect 2087 -3287 2179 -3281
rect 2245 -3247 2337 -3241
rect 2245 -3281 2257 -3247
rect 2325 -3281 2337 -3247
rect 2245 -3287 2337 -3281
rect 2403 -3247 2495 -3241
rect 2403 -3281 2415 -3247
rect 2483 -3281 2495 -3247
rect 2403 -3287 2495 -3281
<< properties >>
string FIXED_BBOX -2662 -3402 2662 3402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 0.5 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
