magic
tech sky130A
magscale 1 2
timestamp 1713239999
<< pwell >>
rect -782 -2202 782 2202
<< psubdiff >>
rect -746 2132 -650 2166
rect 650 2132 746 2166
rect -746 2070 -712 2132
rect 712 2070 746 2132
rect -746 -2132 -712 -2070
rect 712 -2132 746 -2070
rect -746 -2166 -650 -2132
rect 650 -2166 746 -2132
<< psubdiffcont >>
rect -650 2132 650 2166
rect -746 -2070 -712 2070
rect 712 -2070 746 2070
rect -650 -2166 650 -2132
<< xpolycontact >>
rect -616 1604 -546 2036
rect -616 -2036 -546 -1604
rect -450 1604 -380 2036
rect -450 -2036 -380 -1604
rect -284 1604 -214 2036
rect -284 -2036 -214 -1604
rect -118 1604 -48 2036
rect -118 -2036 -48 -1604
rect 48 1604 118 2036
rect 48 -2036 118 -1604
rect 214 1604 284 2036
rect 214 -2036 284 -1604
rect 380 1604 450 2036
rect 380 -2036 450 -1604
rect 546 1604 616 2036
rect 546 -2036 616 -1604
<< xpolyres >>
rect -616 -1604 -546 1604
rect -450 -1604 -380 1604
rect -284 -1604 -214 1604
rect -118 -1604 -48 1604
rect 48 -1604 118 1604
rect 214 -1604 284 1604
rect 380 -1604 450 1604
rect 546 -1604 616 1604
<< locali >>
rect -746 2132 -650 2166
rect 650 2132 746 2166
rect -746 2070 -712 2132
rect 712 2070 746 2132
rect -746 -2132 -712 -2070
rect 712 -2132 746 -2070
rect -746 -2166 -650 -2132
rect 650 -2166 746 -2132
<< viali >>
rect -600 1621 -562 2018
rect -434 1621 -396 2018
rect -268 1621 -230 2018
rect -102 1621 -64 2018
rect 64 1621 102 2018
rect 230 1621 268 2018
rect 396 1621 434 2018
rect 562 1621 600 2018
rect -600 -2018 -562 -1621
rect -434 -2018 -396 -1621
rect -268 -2018 -230 -1621
rect -102 -2018 -64 -1621
rect 64 -2018 102 -1621
rect 230 -2018 268 -1621
rect 396 -2018 434 -1621
rect 562 -2018 600 -1621
<< metal1 >>
rect -606 2018 -556 2030
rect -606 1621 -600 2018
rect -562 1621 -556 2018
rect -606 1609 -556 1621
rect -440 2018 -390 2030
rect -440 1621 -434 2018
rect -396 1621 -390 2018
rect -440 1609 -390 1621
rect -274 2018 -224 2030
rect -274 1621 -268 2018
rect -230 1621 -224 2018
rect -274 1609 -224 1621
rect -108 2018 -58 2030
rect -108 1621 -102 2018
rect -64 1621 -58 2018
rect -108 1609 -58 1621
rect 58 2018 108 2030
rect 58 1621 64 2018
rect 102 1621 108 2018
rect 58 1609 108 1621
rect 224 2018 274 2030
rect 224 1621 230 2018
rect 268 1621 274 2018
rect 224 1609 274 1621
rect 390 2018 440 2030
rect 390 1621 396 2018
rect 434 1621 440 2018
rect 390 1609 440 1621
rect 556 2018 606 2030
rect 556 1621 562 2018
rect 600 1621 606 2018
rect 556 1609 606 1621
rect -606 -1621 -556 -1609
rect -606 -2018 -600 -1621
rect -562 -2018 -556 -1621
rect -606 -2030 -556 -2018
rect -440 -1621 -390 -1609
rect -440 -2018 -434 -1621
rect -396 -2018 -390 -1621
rect -440 -2030 -390 -2018
rect -274 -1621 -224 -1609
rect -274 -2018 -268 -1621
rect -230 -2018 -224 -1621
rect -274 -2030 -224 -2018
rect -108 -1621 -58 -1609
rect -108 -2018 -102 -1621
rect -64 -2018 -58 -1621
rect -108 -2030 -58 -2018
rect 58 -1621 108 -1609
rect 58 -2018 64 -1621
rect 102 -2018 108 -1621
rect 58 -2030 108 -2018
rect 224 -1621 274 -1609
rect 224 -2018 230 -1621
rect 268 -2018 274 -1621
rect 224 -2030 274 -2018
rect 390 -1621 440 -1609
rect 390 -2018 396 -1621
rect 434 -2018 440 -1621
rect 390 -2030 440 -2018
rect 556 -1621 606 -1609
rect 556 -2018 562 -1621
rect 600 -2018 606 -1621
rect 556 -2030 606 -2018
<< properties >>
string FIXED_BBOX -729 -2149 729 2149
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 16.2 m 1 nx 8 wmin 0.350 lmin 0.50 rho 2000 val 93.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
