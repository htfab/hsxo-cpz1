magic
tech sky130A
timestamp 1712933332
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
rect 0 -1800 100 -1700
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC1
timestamp 1712933332
transform 1 0 843 0 1 -5180
box -843 -4980 843 4980
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 XOUT
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 XIN
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 ENA
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 STDBY
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 DOUT
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 AVDD
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 DVDD
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 128 0 0 0 AVSS
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 128 0 0 0 DVSS
port 8 nsew
flabel metal1 0 -1800 100 -1700 0 FreeSans 128 0 0 0 IBIAS
port 9 nsew
<< end >>
