magic
tech sky130A
magscale 1 2
timestamp 1713241921
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
<< nwell >>
rect -226 -319 226 319
<< pmos >>
rect -30 -100 30 100
<< pdiff >>
rect -88 88 -30 100
rect -88 -88 -76 88
rect -42 -88 -30 88
rect -88 -100 -30 -88
rect 30 88 88 100
rect 30 -88 42 88
rect 76 -88 88 88
rect 30 -100 88 -88
<< pdiffc >>
rect -76 -88 -42 88
rect 42 -88 76 88
<< nsubdiff >>
rect -190 249 -94 283
rect 94 249 190 283
rect -190 187 -156 249
rect 156 187 190 249
rect -190 -249 -156 -187
rect 156 -249 190 -187
rect -190 -283 -94 -249
rect 94 -283 190 -249
<< nsubdiffcont >>
rect -94 249 94 283
rect -190 -187 -156 187
rect 156 -187 190 187
rect -94 -283 94 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -30 100 30 131
rect -30 -131 30 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -190 249 -94 283
rect 94 249 190 283
rect -190 187 -156 249
rect 156 187 190 249
rect -33 147 -17 181
rect 17 147 33 181
rect -76 88 -42 104
rect -76 -104 -42 -88
rect 42 88 76 104
rect 42 -104 76 -88
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -190 -249 -156 -187
rect 156 -249 190 -187
rect -190 -283 -94 -249
rect 94 -283 190 -249
<< viali >>
rect -17 147 17 181
rect -76 -88 -42 88
rect 42 -88 76 88
rect -17 -181 17 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -82 88 -36 100
rect -82 -88 -76 88
rect -42 -88 -36 88
rect -82 -100 -36 -88
rect 36 88 82 100
rect 36 -88 42 88
rect 76 -88 82 88
rect 36 -100 82 -88
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
<< properties >>
string FIXED_BBOX -173 -266 173 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
