magic
tech sky130A
magscale 1 2
timestamp 1713252812
<< nwell >>
rect 400 1410 4570 1420
rect 400 620 1120 1410
rect 2340 620 3340 1410
rect 4560 620 4570 1410
rect 400 -1860 980 620
rect 400 -2870 4830 -1860
<< pwell >>
rect 1700 -150 1760 570
rect 2320 -150 3360 570
rect 3930 -150 3980 570
rect 4540 -150 5310 570
rect 1290 -3700 2410 -3570
rect 1290 -4070 1630 -3700
rect 1970 -4044 1990 -4040
rect 1970 -4064 1992 -4044
rect 2000 -4070 2410 -3700
rect 1290 -4200 2410 -4070
rect 3440 -4250 3810 -3350
rect 4840 -4260 5310 -150
<< locali >>
rect 1630 1724 1830 1730
rect 1630 1536 1636 1724
rect 1824 1536 1830 1724
rect 1630 1356 1830 1536
rect 3850 1724 4050 1730
rect 3850 1536 3856 1724
rect 4044 1536 4050 1724
rect 3850 1356 4050 1536
rect 1184 1350 2282 1356
rect 3404 1350 4502 1356
rect 1178 1282 2288 1350
rect 1178 752 1252 1282
rect 1604 1150 1862 1282
rect 1604 752 1678 1150
rect 1178 684 1678 752
rect 1788 752 1862 1150
rect 2214 752 2288 1282
rect 1788 684 2288 752
rect 3398 1282 4508 1350
rect 3398 752 3472 1282
rect 3824 1150 4082 1282
rect 3824 752 3898 1150
rect 3398 684 3898 752
rect 4008 752 4082 1150
rect 4434 752 4508 1282
rect 4008 684 4508 752
rect 1184 678 1672 684
rect 1794 678 2282 684
rect 3404 678 3892 684
rect 4014 678 4502 684
rect 1184 534 1672 538
rect 1794 534 2282 538
rect 1184 532 1636 534
rect 1178 464 1636 532
rect 1178 -48 1252 464
rect 1604 346 1636 464
rect 1824 532 2282 534
rect 3404 532 3892 538
rect 4014 532 4502 538
rect 1824 464 2288 532
rect 1824 346 1862 464
rect 1604 -48 1678 346
rect 1178 -116 1678 -48
rect 1788 -48 1862 346
rect 2214 -48 2288 464
rect 1788 -116 2288 -48
rect 3398 464 3898 532
rect 3398 -48 3472 464
rect 3824 80 3898 464
rect 4008 464 4508 532
rect 4008 80 4082 464
rect 3824 -48 4082 80
rect 4434 -48 4508 464
rect 3398 -116 4508 -48
rect 1184 -122 1672 -116
rect 1794 -122 2282 -116
rect 3404 -122 4502 -116
rect 3850 -426 4050 -122
rect 3850 -614 3856 -426
rect 4044 -614 4050 -426
rect 3850 -620 4050 -614
rect 2760 -1536 2960 -1530
rect 2760 -1724 2766 -1536
rect 2954 -1724 2960 -1536
rect 1958 -1924 2482 -1920
rect 2760 -1924 2960 -1724
rect 3370 -1924 3840 -1920
rect 1054 -1930 4766 -1924
rect 1048 -1998 4772 -1930
rect 1048 -2728 1122 -1998
rect 1948 -2125 2502 -1998
rect 1948 -2728 2022 -2125
rect 1048 -2733 2022 -2728
rect 934 -2796 2022 -2733
rect 2428 -2728 2502 -2125
rect 3328 -2120 3872 -1998
rect 3328 -2728 3402 -2120
rect 2428 -2796 3402 -2728
rect 3798 -2728 3872 -2120
rect 4698 -2728 4772 -1998
rect 3798 -2796 4772 -2728
rect 934 -2802 2016 -2796
rect 2434 -2802 3396 -2796
rect 3804 -2802 4766 -2796
rect 934 -2807 1137 -2802
rect 934 -2879 1008 -2807
rect 934 -2941 940 -2879
rect 1002 -2941 1008 -2879
rect 934 -2947 1008 -2941
rect 2444 -3378 3406 -3372
rect 3844 -3378 4806 -3372
rect 2438 -3446 3412 -3378
rect 616 -3610 1337 -3533
rect 616 -4170 693 -3610
rect 810 -3728 934 -3722
rect 804 -3774 934 -3728
rect 1008 -3728 1132 -3722
rect 1008 -3774 1138 -3728
rect 804 -3796 1138 -3774
rect 804 -3982 878 -3796
rect 1064 -3982 1138 -3796
rect 804 -4050 1138 -3982
rect 810 -4056 1132 -4050
rect 1262 -4170 1337 -3610
rect 1633 -3711 1987 -3710
rect 1633 -3784 1992 -3711
rect 1634 -3990 1712 -3784
rect 1914 -3990 1992 -3784
rect 1633 -4064 1992 -3990
rect 616 -4171 1337 -4170
rect 693 -4237 1337 -4171
rect 2438 -4158 2512 -3446
rect 3338 -4035 3412 -3446
rect 3838 -3446 4812 -3378
rect 3838 -4035 3912 -3446
rect 3338 -4158 3912 -4035
rect 4738 -4158 4812 -3446
rect 2438 -4200 4812 -4158
rect 1920 -4206 4812 -4200
rect 693 -4244 1270 -4237
rect 1920 -4394 1926 -4206
rect 2114 -4226 4812 -4206
rect 2114 -4232 4806 -4226
rect 2114 -4394 2490 -4232
rect 3360 -4240 3892 -4232
rect 1920 -4400 2490 -4394
<< viali >>
rect 1636 1536 1824 1724
rect 3856 1536 4044 1724
rect 1636 346 1824 534
rect 3856 -614 4044 -426
rect 2766 -1724 2954 -1536
rect 940 -2941 1002 -2879
rect 934 -3774 1008 -3700
rect 616 -4248 693 -4171
rect 1926 -4394 2114 -4206
<< metal1 >>
rect 1630 1730 1830 1736
rect 2760 1730 2960 1736
rect 3850 1730 4050 1736
rect 324 1530 330 1730
rect 530 1530 536 1730
rect 1624 1530 1630 1730
rect 1830 1530 1836 1730
rect 3844 1530 3850 1730
rect 4050 1530 4056 1730
rect 330 -3580 530 1530
rect 1630 1524 1830 1530
rect 722 527 728 732
rect 933 527 939 732
rect 728 -1528 933 527
rect 1624 340 1630 540
rect 1830 340 1836 540
rect 2300 530 2330 730
rect 2530 530 2600 730
rect 1934 -260 1940 -60
rect 2140 -260 2146 -60
rect 1940 -420 2140 -260
rect 1104 -620 1110 -420
rect 1310 -620 2140 -420
rect 728 -1739 933 -1733
rect 2400 -1920 2600 530
rect 2760 -1530 2960 1530
rect 3850 1524 4050 1530
rect 3118 730 3303 732
rect 4710 730 4910 736
rect 3118 530 3160 730
rect 3360 530 3390 730
rect 4705 530 4710 702
rect 3118 -1528 3323 530
rect 3544 -260 3550 -60
rect 3750 -260 3756 -60
rect 4154 -260 4160 -60
rect 4360 -260 4366 -60
rect 3550 -790 3750 -260
rect 3850 -420 4050 -414
rect 3850 -626 4050 -620
rect 3544 -990 3550 -790
rect 3750 -990 3756 -790
rect 4160 -1140 4360 -260
rect 4160 -1346 4360 -1340
rect 2760 -1736 2960 -1730
rect 3112 -1733 3118 -1528
rect 3323 -1733 3329 -1528
rect 4705 -1920 4910 530
rect 5550 -420 5750 -414
rect 910 -2125 3540 -1920
rect 910 -2605 1115 -2125
rect 1192 -2175 1246 -2165
rect 1192 -2329 1246 -2319
rect 1508 -2175 1562 -2165
rect 1508 -2329 1562 -2319
rect 1824 -2175 1878 -2165
rect 1824 -2329 1878 -2319
rect 1350 -2407 1404 -2397
rect 1350 -2561 1404 -2551
rect 1666 -2407 1720 -2397
rect 1666 -2561 1720 -2551
rect 1955 -2605 2160 -2125
rect 910 -2810 2160 -2605
rect 2290 -2605 2495 -2125
rect 2572 -2175 2626 -2165
rect 2572 -2329 2626 -2319
rect 2888 -2175 2942 -2165
rect 2888 -2329 2942 -2319
rect 3204 -2175 3258 -2165
rect 3204 -2329 3258 -2319
rect 2730 -2407 2784 -2397
rect 2730 -2561 2784 -2551
rect 3046 -2407 3100 -2397
rect 3046 -2561 3100 -2551
rect 3335 -2605 3540 -2125
rect 2290 -2810 3540 -2605
rect 3660 -2125 4910 -1920
rect 3660 -2605 3865 -2125
rect 3942 -2175 3996 -2165
rect 3942 -2329 3996 -2319
rect 4258 -2175 4312 -2165
rect 4258 -2329 4312 -2319
rect 4574 -2175 4628 -2165
rect 4574 -2329 4628 -2319
rect 4100 -2407 4154 -2397
rect 4100 -2561 4154 -2551
rect 4416 -2407 4470 -2397
rect 4416 -2561 4470 -2551
rect 4705 -2605 4910 -2125
rect 3660 -2810 4910 -2605
rect 5137 -1528 5342 -1522
rect 928 -2879 1014 -2873
rect 928 -2941 940 -2879
rect 1002 -2941 1014 -2879
rect 928 -2947 1014 -2941
rect 330 -3780 860 -3580
rect 934 -3694 1008 -2947
rect 2112 -3443 2118 -3238
rect 2323 -3360 2495 -3238
rect 5137 -3360 5342 -1733
rect 2323 -3443 3540 -3360
rect 2290 -3565 3540 -3443
rect 922 -3700 1020 -3694
rect 922 -3774 934 -3700
rect 1008 -3774 1020 -3700
rect 922 -3780 1020 -3774
rect 660 -4000 860 -3780
rect 900 -3830 1040 -3820
rect 900 -3950 910 -3830
rect 1030 -3950 1040 -3830
rect 900 -3960 1040 -3950
rect 1080 -3852 1280 -3580
rect 1500 -3780 2120 -3580
rect 1080 -4000 1338 -3852
rect 660 -4159 1338 -4000
rect 610 -4171 1338 -4159
rect 610 -4248 616 -4171
rect 693 -4247 1338 -4171
rect 1500 -4000 1700 -3780
rect 1740 -3830 1880 -3820
rect 1740 -3950 1750 -3830
rect 1870 -3950 1880 -3830
rect 1740 -3960 1880 -3950
rect 1920 -4000 2120 -3780
rect 1500 -4200 2120 -4000
rect 2290 -4035 2490 -3565
rect 2582 -3614 2636 -3604
rect 2582 -3768 2636 -3758
rect 2898 -3614 2952 -3604
rect 2898 -3768 2952 -3758
rect 3214 -3614 3268 -3604
rect 3214 -3768 3268 -3758
rect 2740 -3846 2794 -3836
rect 2740 -4000 2794 -3990
rect 3056 -3846 3110 -3836
rect 3056 -4000 3110 -3990
rect 3340 -4035 3540 -3565
rect 693 -4248 699 -4247
rect 610 -4260 699 -4248
rect 1914 -4400 1920 -4200
rect 2120 -4400 2126 -4200
rect 2290 -4240 3540 -4035
rect 3670 -3565 5342 -3360
rect 3670 -4035 3870 -3565
rect 3982 -3614 4036 -3604
rect 3982 -3768 4036 -3758
rect 4298 -3614 4352 -3604
rect 4298 -3768 4352 -3758
rect 4614 -3614 4668 -3604
rect 4614 -3768 4668 -3758
rect 4140 -3846 4194 -3836
rect 4140 -4000 4194 -3990
rect 4456 -3846 4510 -3836
rect 4456 -4000 4510 -3990
rect 4700 -4035 4900 -3565
rect 3670 -4240 4900 -4035
rect 5550 -4030 5750 -620
rect 5550 -4236 5750 -4230
rect 1920 -4406 2120 -4400
<< via1 >>
rect 330 1530 530 1730
rect 1630 1724 1830 1730
rect 1630 1536 1636 1724
rect 1636 1536 1824 1724
rect 1824 1536 1830 1724
rect 1630 1530 1830 1536
rect 2760 1530 2960 1730
rect 3850 1724 4050 1730
rect 3850 1536 3856 1724
rect 3856 1536 4044 1724
rect 4044 1536 4050 1724
rect 3850 1530 4050 1536
rect 728 527 933 732
rect 1630 534 1830 540
rect 1630 346 1636 534
rect 1636 346 1824 534
rect 1824 346 1830 534
rect 1630 340 1830 346
rect 2330 530 2530 730
rect 1940 -260 2140 -60
rect 1110 -620 1310 -420
rect 728 -1733 933 -1528
rect 3160 530 3360 730
rect 4710 530 4910 730
rect 3550 -260 3750 -60
rect 4160 -260 4360 -60
rect 3850 -426 4050 -420
rect 3850 -614 3856 -426
rect 3856 -614 4044 -426
rect 4044 -614 4050 -426
rect 3850 -620 4050 -614
rect 3550 -990 3750 -790
rect 4160 -1340 4360 -1140
rect 2760 -1536 2960 -1530
rect 2760 -1724 2766 -1536
rect 2766 -1724 2954 -1536
rect 2954 -1724 2960 -1536
rect 2760 -1730 2960 -1724
rect 3118 -1733 3323 -1528
rect 5550 -620 5750 -420
rect 1192 -2319 1246 -2175
rect 1508 -2319 1562 -2175
rect 1824 -2319 1878 -2175
rect 1350 -2551 1404 -2407
rect 1666 -2551 1720 -2407
rect 2572 -2319 2626 -2175
rect 2888 -2319 2942 -2175
rect 3204 -2319 3258 -2175
rect 2730 -2551 2784 -2407
rect 3046 -2551 3100 -2407
rect 3942 -2319 3996 -2175
rect 4258 -2319 4312 -2175
rect 4574 -2319 4628 -2175
rect 4100 -2551 4154 -2407
rect 4416 -2551 4470 -2407
rect 5137 -1733 5342 -1528
rect 2118 -3443 2323 -3238
rect 910 -3950 1030 -3830
rect 1750 -3950 1870 -3830
rect 2582 -3758 2636 -3614
rect 2898 -3758 2952 -3614
rect 3214 -3758 3268 -3614
rect 2740 -3990 2794 -3846
rect 3056 -3990 3110 -3846
rect 1920 -4206 2120 -4200
rect 1920 -4394 1926 -4206
rect 1926 -4394 2114 -4206
rect 2114 -4394 2120 -4206
rect 1920 -4400 2120 -4394
rect 3982 -3758 4036 -3614
rect 4298 -3758 4352 -3614
rect 4614 -3758 4668 -3614
rect 4140 -3990 4194 -3846
rect 4456 -3990 4510 -3846
rect 5550 -4230 5750 -4030
<< metal2 >>
rect 330 1730 530 1736
rect 130 1530 330 1730
rect 530 1530 1630 1730
rect 1830 1530 2760 1730
rect 2960 1530 3850 1730
rect 4050 1530 4056 1730
rect 330 1524 530 1530
rect 1630 1300 1830 1530
rect 3850 1300 4050 1530
rect 728 732 933 738
rect 933 527 1172 732
rect 2330 730 2530 736
rect 1630 540 1830 546
rect 728 521 933 527
rect 2250 530 2330 730
rect 2330 524 2530 530
rect 3160 730 3360 736
rect 3360 530 3440 730
rect 4470 530 4710 730
rect 4910 530 4916 730
rect 3160 524 3360 530
rect 130 -260 1530 -60
rect 1110 -420 1310 -414
rect 130 -620 1110 -420
rect 1630 -420 1830 340
rect 1940 -60 2140 -54
rect 1940 -266 2140 -260
rect 3550 -60 3750 -54
rect 4160 -60 4360 -54
rect 3550 -266 3750 -260
rect 3850 -420 4050 -60
rect 4160 -266 4360 -260
rect 1630 -620 3850 -420
rect 4050 -620 5550 -420
rect 5750 -620 5756 -420
rect 1110 -626 1310 -620
rect 3550 -790 3750 -784
rect 130 -990 3550 -790
rect 3550 -996 3750 -990
rect 130 -1340 4160 -1140
rect 4360 -1340 4366 -1140
rect 3118 -1528 3323 -1522
rect 722 -1733 728 -1528
rect 933 -1733 2323 -1528
rect 130 -2175 1890 -2130
rect 130 -2319 1192 -2175
rect 1246 -2319 1508 -2175
rect 1562 -2319 1824 -2175
rect 1878 -2319 1890 -2175
rect 130 -2330 1890 -2319
rect 1170 -2407 1890 -2400
rect 1170 -2530 1350 -2407
rect 130 -2551 1350 -2530
rect 1404 -2551 1666 -2407
rect 1720 -2551 1890 -2407
rect 130 -2600 1890 -2551
rect 130 -2730 1370 -2600
rect 2118 -3238 2323 -1733
rect 2600 -1730 2760 -1530
rect 2960 -1730 2966 -1530
rect 2600 -2130 2800 -1730
rect 3323 -1733 5137 -1528
rect 5342 -1733 5348 -1528
rect 3118 -1739 3323 -1733
rect 2560 -2175 4640 -2130
rect 2560 -2319 2572 -2175
rect 2626 -2319 2888 -2175
rect 2942 -2319 3204 -2175
rect 3258 -2319 3942 -2175
rect 3996 -2319 4258 -2175
rect 4312 -2319 4574 -2175
rect 4628 -2319 4640 -2175
rect 2560 -2330 4640 -2319
rect 2560 -2407 3280 -2400
rect 2560 -2551 2730 -2407
rect 2784 -2551 3046 -2407
rect 3100 -2551 3280 -2407
rect 2560 -2600 3280 -2551
rect 3930 -2407 5950 -2400
rect 3930 -2551 4100 -2407
rect 4154 -2551 4416 -2407
rect 4470 -2551 5950 -2407
rect 3930 -2600 5950 -2551
rect 3080 -2760 3280 -2600
rect 3080 -2960 5950 -2760
rect 2118 -3449 2323 -3443
rect 3080 -3380 5950 -3180
rect 3080 -3570 3280 -3380
rect 2570 -3614 3280 -3570
rect 2570 -3758 2582 -3614
rect 2636 -3758 2898 -3614
rect 2952 -3758 3214 -3614
rect 3268 -3758 3280 -3614
rect 2570 -3770 3280 -3758
rect 3970 -3614 5950 -3570
rect 3970 -3758 3982 -3614
rect 4036 -3758 4298 -3614
rect 4352 -3758 4614 -3614
rect 4668 -3758 5950 -3614
rect 3970 -3770 5950 -3758
rect 871 -3790 1071 -3789
rect 130 -3830 1910 -3790
rect 130 -3950 910 -3830
rect 1030 -3950 1750 -3830
rect 1870 -3950 1910 -3830
rect 130 -3990 1910 -3950
rect 2570 -3846 4690 -3840
rect 2570 -3990 2740 -3846
rect 2794 -3990 3056 -3846
rect 3110 -3990 4140 -3846
rect 4194 -3990 4456 -3846
rect 4510 -3990 4690 -3846
rect 2570 -4030 4690 -3990
rect 2570 -4040 5550 -4030
rect 1920 -4200 2120 -4194
rect 2570 -4200 2770 -4040
rect 130 -4400 1920 -4200
rect 2120 -4400 2770 -4200
rect 4490 -4230 5550 -4040
rect 5750 -4230 5756 -4030
rect 1920 -4406 2120 -4400
use p_diode  D1
timestamp 1713252812
transform 1 0 971 0 1 -3889
box -371 -370 381 369
use n_diode  D2
timestamp 1713252812
transform 1 0 1813 0 1 -3887
box -193 -193 193 193
use level_shifter_ad  level_shifter_ad_0
timestamp 1713252812
transform 1 0 140 0 1 1710
box 880 -1970 2310 -210
use level_shifter_ad  level_shifter_ad_1
timestamp 1713252812
transform 1 0 2360 0 1 1710
box 880 -1970 2310 -210
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM1
timestamp 1713252812
transform 1 0 4285 0 1 -2363
box -545 -497 545 497
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM2
timestamp 1713252812
transform 1 0 1535 0 1 -2363
box -545 -497 545 497
use sky130_fd_pr__nfet_g5v0d10v5_F7BQJ6  XM3
timestamp 1713252812
transform 1 0 4325 0 1 -3802
box -515 -458 515 458
use sky130_fd_pr__nfet_g5v0d10v5_F7BQJ6  XM21
timestamp 1713252812
transform 1 0 2925 0 1 -3802
box -515 -458 515 458
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM25
timestamp 1713252812
transform 1 0 2915 0 1 -2363
box -545 -497 545 497
<< labels >>
flabel metal2 130 1530 330 1730 0 FreeSans 256 0 0 0 AVDD
port 5 nsew
flabel metal2 130 -260 330 -60 0 FreeSans 256 0 0 0 ENA
port 8 nsew
flabel metal2 130 -620 330 -420 0 FreeSans 256 0 0 0 ENA_B
port 8 nsew
flabel metal2 130 -990 330 -790 0 FreeSans 256 0 0 0 STDBY
port 11 nsew
flabel metal2 130 -1340 330 -1140 0 FreeSans 256 0 0 0 STDBY_B
port 11 nsew
flabel metal2 130 -2330 330 -2130 0 FreeSans 256 0 0 0 IBIAS
port 6 nsew
flabel metal2 130 -2730 330 -2530 0 FreeSans 256 0 0 0 EG_IBIAS
port 3 nsew
flabel metal2 130 -4400 330 -4200 0 FreeSans 256 0 0 0 AVSS
port 13 nsew
flabel metal2 5750 -2600 5950 -2400 0 FreeSans 256 0 0 0 SG_AVDD
port 1 nsew
flabel metal2 5750 -2960 5950 -2760 0 FreeSans 256 0 0 0 EG_AVDD
port 7 nsew
flabel metal2 5750 -3380 5950 -3180 0 FreeSans 256 0 0 0 EG_AVSS
port 12 nsew
flabel metal2 5750 -3770 5950 -3570 0 FreeSans 256 0 0 0 SG_AVSS
port 10 nsew
flabel metal2 130 -3990 330 -3790 0 FreeSans 256 0 0 0 XIN
port 3 nsew
<< end >>
