magic
tech sky130A
magscale 1 2
timestamp 1713795963
<< nwell >>
rect 1800 -3220 2270 -1720
rect 2690 -2360 4324 -1720
rect 1800 -4450 2100 -3220
<< pwell >>
rect 2700 -2980 4324 -2360
rect 3854 -3550 4744 -2980
rect 3854 -4620 4740 -3550
rect 3854 -5110 4960 -4620
rect 3204 -6330 3854 -5110
rect 4910 -5120 4960 -5110
rect 4950 -6330 4960 -5120
<< locali >>
rect 2292 -1744 2670 -1738
rect 4346 -1744 4724 -1738
rect 2286 -1812 2676 -1744
rect 2286 -1940 2360 -1812
rect 1710 -2140 2360 -1940
rect 2286 -2270 2360 -2140
rect 2602 -2270 2676 -1812
rect 4340 -1812 4730 -1744
rect 4340 -1940 4414 -1812
rect 3960 -2140 4414 -1940
rect 2286 -2338 2676 -2270
rect 4340 -2270 4414 -2140
rect 4656 -2270 4730 -1812
rect 4340 -2338 4730 -2270
rect 2292 -2340 2670 -2338
rect 4346 -2340 4724 -2338
rect 2292 -2382 2670 -2380
rect 4346 -2382 4724 -2380
rect 2286 -2450 2676 -2382
rect 2286 -2890 2360 -2450
rect 2602 -2890 2676 -2450
rect 4340 -2450 4730 -2382
rect 4340 -2760 4414 -2450
rect 2286 -2958 2676 -2890
rect 4164 -2890 4414 -2760
rect 4656 -2890 4730 -2450
rect 4164 -2958 4730 -2890
rect 2292 -2964 2670 -2958
rect 4164 -2964 4724 -2958
rect 4164 -3026 4364 -2964
rect 4164 -3214 4170 -3026
rect 4358 -3214 4364 -3026
rect 4164 -3220 4364 -3214
rect 2122 -3234 3180 -3228
rect 2116 -3302 3186 -3234
rect 2116 -4360 2190 -3302
rect 3112 -3390 3186 -3302
rect 3112 -3396 3960 -3390
rect 3112 -3784 3566 -3396
rect 3954 -3784 3960 -3396
rect 3112 -3790 3960 -3784
rect 3112 -4360 3186 -3790
rect 2116 -4428 3186 -4360
rect 2122 -4434 3180 -4428
rect 2124 -5132 3182 -5126
rect 3876 -5132 4934 -5126
rect 2118 -5200 3188 -5132
rect 2118 -6240 2192 -5200
rect 3114 -5760 3188 -5200
rect 3870 -5200 4940 -5132
rect 3870 -5760 3944 -5200
rect 3114 -6160 3944 -5760
rect 3114 -6240 3188 -6160
rect 2118 -6308 3188 -6240
rect 3870 -6240 3944 -6160
rect 4866 -5759 4940 -5200
rect 4866 -5765 5760 -5759
rect 4866 -6155 5364 -5765
rect 5754 -6155 5760 -5765
rect 4866 -6161 5760 -6155
rect 4866 -6240 4940 -6161
rect 3870 -6308 4940 -6240
rect 2124 -6314 3182 -6308
rect 3876 -6314 4934 -6308
<< viali >>
rect 1510 -2140 1710 -1940
rect 3760 -2140 3960 -1940
rect 4170 -3214 4358 -3026
rect 3566 -3784 3954 -3396
rect 5364 -6155 5754 -5765
<< metal1 >>
rect 1504 -1930 1716 -1928
rect 1310 -1940 1716 -1930
rect 3748 -1940 3972 -1934
rect 1310 -2140 1510 -1940
rect 1710 -2140 1716 -1940
rect 1310 -2152 1716 -2140
rect 3560 -2140 3750 -1940
rect 3960 -2140 3972 -1940
rect 3560 -2146 3972 -2140
rect 1310 -3390 1710 -2152
rect 3188 -2460 3194 -2260
rect 3394 -2460 3400 -2260
rect 3194 -3190 3394 -2460
rect 1900 -3390 3394 -3190
rect 3560 -3390 3960 -2146
rect 4910 -2260 5110 -2254
rect 4910 -3020 5110 -2460
rect 4158 -3220 4164 -3020
rect 4364 -3220 4370 -3020
rect 4560 -3220 5110 -3020
rect 1304 -3790 1310 -3390
rect 1710 -3790 1716 -3390
rect 1900 -4270 2100 -3390
rect 2240 -3443 2294 -3433
rect 2240 -3597 2294 -3587
rect 2432 -3443 2486 -3433
rect 2432 -3597 2486 -3587
rect 2624 -3443 2678 -3433
rect 2624 -3597 2678 -3587
rect 2816 -3443 2870 -3433
rect 2816 -3597 2870 -3587
rect 3008 -3443 3062 -3433
rect 3008 -3597 3062 -3587
rect 2336 -4075 2390 -4065
rect 2336 -4229 2390 -4219
rect 2528 -4075 2582 -4065
rect 2528 -4229 2582 -4219
rect 2720 -4075 2774 -4065
rect 2720 -4229 2774 -4219
rect 2912 -4075 2966 -4065
rect 2912 -4229 2966 -4219
rect 3194 -4270 3394 -3390
rect 3554 -3790 3560 -3390
rect 3960 -3790 3966 -3390
rect 4154 -3850 4160 -3650
rect 4360 -3850 4366 -3650
rect 4160 -4270 4360 -3850
rect 1900 -4470 4360 -4270
rect 4560 -4690 4760 -3220
rect 5352 -3421 5358 -3019
rect 5760 -3421 5766 -3019
rect 3196 -4890 4760 -4690
rect 4960 -3650 5160 -3644
rect 3196 -5090 3396 -4890
rect 4960 -5090 5160 -3850
rect 1902 -5290 3396 -5090
rect 1902 -6160 2102 -5290
rect 2242 -5332 2296 -5322
rect 2242 -5486 2296 -5476
rect 2434 -5332 2488 -5322
rect 2434 -5486 2488 -5476
rect 2626 -5332 2680 -5322
rect 2626 -5486 2680 -5476
rect 2818 -5332 2872 -5322
rect 2818 -5486 2872 -5476
rect 3010 -5332 3064 -5322
rect 3010 -5486 3064 -5476
rect 2338 -5964 2392 -5954
rect 2338 -6118 2392 -6108
rect 2530 -5964 2584 -5954
rect 2530 -6118 2584 -6108
rect 2722 -5964 2776 -5954
rect 2722 -6118 2776 -6108
rect 2914 -5964 2968 -5954
rect 2914 -6118 2968 -6108
rect 3196 -6160 3396 -5290
rect 1900 -6360 3396 -6160
rect 3654 -5290 5160 -5090
rect 3654 -6150 3854 -5290
rect 3994 -5332 4048 -5322
rect 3994 -5486 4048 -5476
rect 4186 -5332 4240 -5322
rect 4186 -5486 4240 -5476
rect 4378 -5332 4432 -5322
rect 4378 -5486 4432 -5476
rect 4570 -5332 4624 -5322
rect 4570 -5486 4624 -5476
rect 4762 -5332 4816 -5322
rect 4762 -5486 4816 -5476
rect 4958 -5430 5160 -5290
rect 4090 -5964 4144 -5954
rect 4090 -6118 4144 -6108
rect 4282 -5964 4336 -5954
rect 4282 -6118 4336 -6108
rect 4474 -5964 4528 -5954
rect 4474 -6118 4528 -6108
rect 4666 -5964 4720 -5954
rect 4666 -6118 4720 -6108
rect 4958 -6150 5158 -5430
rect 5358 -5759 5760 -3421
rect 3654 -6360 5158 -6150
rect 5352 -5760 5766 -5759
rect 5352 -5960 5360 -5760
rect 5352 -6160 5358 -5960
rect 5760 -6160 5766 -5760
rect 5352 -6161 5766 -6160
rect 5358 -6166 5558 -6161
<< via1 >>
rect 3750 -2140 3760 -1940
rect 3760 -2140 3950 -1940
rect 3194 -2460 3394 -2260
rect 4910 -2460 5110 -2260
rect 4164 -3026 4364 -3020
rect 4164 -3214 4170 -3026
rect 4170 -3214 4358 -3026
rect 4358 -3214 4364 -3026
rect 4164 -3220 4364 -3214
rect 1310 -3790 1710 -3390
rect 2240 -3587 2294 -3443
rect 2432 -3587 2486 -3443
rect 2624 -3587 2678 -3443
rect 2816 -3587 2870 -3443
rect 3008 -3587 3062 -3443
rect 2336 -4219 2390 -4075
rect 2528 -4219 2582 -4075
rect 2720 -4219 2774 -4075
rect 2912 -4219 2966 -4075
rect 3560 -3396 3960 -3390
rect 3560 -3784 3566 -3396
rect 3566 -3784 3954 -3396
rect 3954 -3784 3960 -3396
rect 3560 -3790 3960 -3784
rect 4160 -3850 4360 -3650
rect 5358 -3421 5760 -3019
rect 4960 -3850 5160 -3650
rect 2242 -5476 2296 -5332
rect 2434 -5476 2488 -5332
rect 2626 -5476 2680 -5332
rect 2818 -5476 2872 -5332
rect 3010 -5476 3064 -5332
rect 2338 -6108 2392 -5964
rect 2530 -6108 2584 -5964
rect 2722 -6108 2776 -5964
rect 2914 -6108 2968 -5964
rect 3994 -5476 4048 -5332
rect 4186 -5476 4240 -5332
rect 4378 -5476 4432 -5332
rect 4570 -5476 4624 -5332
rect 4762 -5476 4816 -5332
rect 4090 -6108 4144 -5964
rect 4282 -6108 4336 -5964
rect 4474 -6108 4528 -5964
rect 4666 -6108 4720 -5964
rect 5360 -5765 5760 -5760
rect 5360 -5960 5364 -5765
rect 5358 -6155 5364 -5960
rect 5364 -6155 5754 -5765
rect 5754 -6155 5760 -5765
rect 5358 -6160 5760 -6155
<< metal2 >>
rect 1710 -2260 1910 -1320
rect 2110 -2140 2310 -1940
rect 1710 -2460 2310 -2260
rect 2650 -2460 2850 -1320
rect 3190 -2254 3390 -1320
rect 3750 -1940 3950 -1934
rect 3950 -2140 4354 -1940
rect 3750 -2146 3950 -2140
rect 3190 -2260 3394 -2254
rect 4910 -2260 5110 -1320
rect 3190 -2460 3194 -2260
rect 3394 -2460 4364 -2260
rect 4704 -2460 4910 -2260
rect 5110 -2460 5116 -2260
rect 3194 -2466 3394 -2460
rect 2110 -3020 2310 -2570
rect 3194 -2770 4364 -2570
rect 3194 -3020 3394 -2770
rect 4164 -3019 4364 -2770
rect 5358 -3019 5760 -3013
rect 2110 -3220 3394 -3020
rect 4159 -3020 5358 -3019
rect 4159 -3220 4164 -3020
rect 4364 -3220 5358 -3020
rect 1310 -3390 1710 -3384
rect 3560 -3390 3960 -3384
rect 1710 -3443 3560 -3390
rect 1710 -3587 2240 -3443
rect 2294 -3587 2432 -3443
rect 2486 -3587 2624 -3443
rect 2678 -3587 2816 -3443
rect 2870 -3587 3008 -3443
rect 3062 -3587 3560 -3443
rect 1710 -3790 3560 -3587
rect 4159 -3421 5358 -3220
rect 5358 -3427 5760 -3421
rect 1310 -3796 1710 -3790
rect 3560 -3796 3960 -3790
rect 4160 -3650 4360 -3644
rect 4360 -3850 4960 -3650
rect 5160 -3850 5166 -3650
rect 4160 -3856 4360 -3850
rect 2220 -4075 6360 -4070
rect 2220 -4219 2336 -4075
rect 2390 -4219 2528 -4075
rect 2582 -4219 2720 -4075
rect 2774 -4219 2912 -4075
rect 2966 -4219 6360 -4075
rect 2220 -4470 6360 -4219
rect 2680 -5060 6360 -4660
rect 2680 -5080 3080 -5060
rect 2220 -5332 3080 -5080
rect 2220 -5476 2242 -5332
rect 2296 -5476 2434 -5332
rect 2488 -5476 2626 -5332
rect 2680 -5476 2818 -5332
rect 2872 -5476 3010 -5332
rect 3064 -5476 3080 -5332
rect 2220 -5480 3080 -5476
rect 3984 -5332 6358 -5280
rect 3984 -5476 3994 -5332
rect 4048 -5476 4186 -5332
rect 4240 -5476 4378 -5332
rect 4432 -5476 4570 -5332
rect 4624 -5476 4762 -5332
rect 4816 -5476 6358 -5332
rect 3984 -5480 6358 -5476
rect 5360 -5760 5760 -5754
rect 1310 -5960 5360 -5760
rect 1310 -5964 5358 -5960
rect 1310 -6108 2338 -5964
rect 2392 -6108 2530 -5964
rect 2584 -6108 2722 -5964
rect 2776 -6108 2914 -5964
rect 2968 -6108 4090 -5964
rect 4144 -6108 4282 -5964
rect 4336 -6108 4474 -5964
rect 4528 -6108 4666 -5964
rect 4720 -6108 5358 -5964
rect 1310 -6160 5358 -6108
rect 5360 -6166 5760 -6160
use level_shifter_dd  level_shifter_dd_0
timestamp 1713791489
transform 1 0 1890 0 1 -1070
box 220 -1910 960 -652
use level_shifter_dd  level_shifter_dd_1
timestamp 1713791489
transform 1 0 3944 0 1 -1070
box 220 -1910 960 -652
use sky130_fd_pr__nfet_01v8_HNLS5R  sky130_fd_pr__nfet_01v8_HNLS5R_0
timestamp 1713791489
transform 1 0 4405 0 1 -5720
box -551 -610 551 610
use sky130_fd_pr__pfet_01v8_XGNZDL  sky130_fd_pr__pfet_01v8_XGNZDL_0
timestamp 1713794310
transform 1 0 2651 0 1 -3831
box -551 -619 551 619
use sky130_fd_pr__nfet_01v8_HNLS5R  XM18
timestamp 1713791489
transform 1 0 2653 0 1 -5720
box -551 -610 551 610
<< labels >>
flabel metal2 6158 -5480 6358 -5280 0 FreeSans 256 0 0 0 DOUT
port 8 nsew
flabel metal2 5960 -5060 6360 -4660 0 FreeSans 256 0 0 0 SG_DVSS
port 6 nsew
flabel metal2 2650 -1520 2850 -1320 0 FreeSans 256 0 0 0 ENA_B
port 3 nsew
flabel metal2 1710 -1520 1910 -1320 0 FreeSans 256 0 0 0 ENA
port 2 nsew
flabel metal2 3190 -1520 3390 -1320 0 FreeSans 256 0 0 0 STDBY
port 4 nsew
flabel metal2 4910 -1520 5110 -1320 0 FreeSans 256 0 0 0 STDBY_B
port 5 nsew
flabel metal2 5960 -4470 6360 -4070 0 FreeSans 256 0 0 0 SG_DVDD
port 7 nsew
flabel metal2 1310 -3790 1710 -3390 0 FreeSans 256 0 0 0 DVDD
port 1 nsew
flabel metal2 1310 -6160 1710 -5760 0 FreeSans 256 0 0 0 DVSS
port 0 nsew
<< end >>
