magic
tech sky130A
magscale 1 2
timestamp 1718125978
<< isosubstrate >>
rect 1877 3040 4873 3830
rect 3340 2540 4873 3040
rect 1877 1812 4873 2540
rect 1877 920 3530 1812
rect 1877 -1963 4873 920
<< nwell >>
rect 1591 3830 5159 4119
rect 1591 3793 1880 3830
rect 1591 3040 1877 3793
rect 1591 2540 3340 3040
rect 1591 -1963 1877 2540
rect 4873 1810 5159 3830
rect 4160 1540 5159 1810
rect 4520 920 5159 1540
rect 4873 -1963 5159 920
rect 1591 -2249 5159 -1963
<< psubdiff >>
rect 2416 3180 2440 3380
rect 3240 3180 3264 3380
<< nsubdiff >>
rect 1628 4062 5122 4082
rect 1628 4028 1708 4062
rect 5042 4028 5122 4062
rect 1628 4008 5122 4028
rect 1628 4002 1702 4008
rect 1628 -2132 1648 4002
rect 1682 -2132 1702 4002
rect 5048 4002 5122 4008
rect 2416 2680 2440 2880
rect 3240 2680 3264 2880
rect 1628 -2138 1702 -2132
rect 5048 -2132 5068 4002
rect 5102 -2132 5122 4002
rect 5048 -2138 5122 -2132
rect 1628 -2158 5122 -2138
rect 1628 -2192 1708 -2158
rect 5042 -2192 5122 -2158
rect 1628 -2212 5122 -2192
<< mvpsubdiff >>
rect 4126 4428 4302 4462
<< psubdiffcont >>
rect 2440 3180 3240 3380
<< nsubdiffcont >>
rect 1708 4028 5042 4062
rect 1648 -2132 1682 4002
rect 2440 2680 3240 2880
rect 5068 -2132 5102 4002
rect 1708 -2192 5042 -2158
<< locali >>
rect 1648 4028 1708 4062
rect 5042 4028 5102 4062
rect 1648 4002 1682 4028
rect 5068 4002 5102 4028
rect 3532 3794 4388 3800
rect 3526 3726 4394 3794
rect 3526 3380 3600 3726
rect 2424 3180 2440 3380
rect 3240 3180 3600 3380
rect 2424 2680 2440 2880
rect 3240 2680 3256 2880
rect 3526 2458 3600 3180
rect 1982 2452 3600 2458
rect 1976 2384 3600 2452
rect 1976 -1840 2050 2384
rect 3434 1910 3600 2384
rect 4320 1910 4394 3726
rect 3434 1842 4394 1910
rect 3434 1836 4388 1842
rect 3434 107 3508 1836
rect 3552 1790 4146 1796
rect 3546 1722 4152 1790
rect 3546 1450 3620 1722
rect 4078 1710 4152 1722
rect 4078 1704 4310 1710
rect 4078 1616 4216 1704
rect 4304 1616 4310 1704
rect 4078 1542 4310 1616
rect 4078 1536 4580 1542
rect 4078 1468 4586 1536
rect 4078 1450 4240 1468
rect 3546 1282 4240 1450
rect 3546 1010 3620 1282
rect 4078 1010 4240 1282
rect 4512 1010 4586 1468
rect 3546 942 4587 1010
rect 3552 936 4587 942
rect 3562 890 4577 896
rect 3556 822 4577 890
rect 3556 570 3630 822
rect 4070 570 4250 822
rect 3556 402 4250 570
rect 3556 150 3630 402
rect 4070 390 4250 402
rect 4502 390 4576 822
rect 4070 322 4576 390
rect 4070 316 4570 322
rect 4070 150 4144 316
rect 3556 107 4144 150
rect 3434 50 4144 107
rect 3434 44 4388 50
rect 3434 -24 4394 44
rect 3434 -1840 3600 -24
rect 4320 -1840 4394 -24
rect 1976 -1908 4394 -1840
rect 1982 -1914 4388 -1908
rect 1648 -2158 1682 -2132
rect 5068 -2158 5102 -2132
rect 1648 -2192 1708 -2158
rect 5042 -2192 5102 -2158
<< viali >>
rect 2786 3236 2874 3324
rect 2776 2736 2864 2824
rect 4216 1616 4304 1704
<< metal1 >>
rect 2774 3324 3470 3330
rect 2774 3236 2786 3324
rect 2874 3236 3470 3324
rect 2774 3230 3470 3236
rect 3370 3090 3470 3230
rect 3670 3180 3920 3620
rect 4000 3180 4250 3620
rect 3370 2990 4630 3090
rect 2770 2830 2870 2836
rect 2764 2730 2770 2830
rect 2870 2730 2876 2830
rect 2770 2724 2870 2730
rect 3500 2310 3750 2420
rect 2100 970 2200 2310
rect 2280 1870 2530 2310
rect 2620 1870 2870 2310
rect 2950 1870 3200 2310
rect 3280 1980 3750 2310
rect 3830 1980 4080 2420
rect 4170 2079 4420 2420
rect 4170 1980 4321 2079
rect 2100 864 2200 870
rect 3280 -100 3380 1980
rect 4321 1974 4420 1980
rect 3799 1826 3899 1830
rect 3799 1820 3900 1826
rect 3799 1630 3900 1720
rect 3799 1620 3899 1630
rect 3823 1619 3875 1620
rect 3653 1560 3659 1612
rect 3711 1560 3717 1612
rect 3981 1560 3987 1612
rect 4039 1560 4045 1612
rect 4204 1610 4210 1710
rect 4310 1610 4316 1710
rect 3823 1550 3875 1553
rect 3799 1310 3899 1550
rect 4350 1429 4402 1435
rect 4350 1371 4402 1377
rect 4530 1310 4630 2990
rect 3799 1210 4320 1310
rect 4430 1210 4530 1310
rect 4630 1210 4636 1310
rect 3799 1180 3899 1210
rect 3823 1179 3875 1180
rect 3653 1120 3659 1172
rect 3711 1120 3717 1172
rect 3981 1120 3987 1172
rect 4039 1120 4045 1172
rect 3824 1113 3876 1116
rect 3823 1110 3876 1113
rect 3799 970 3899 1110
rect 4320 1010 4326 1110
rect 4426 1010 4432 1110
rect 4326 970 4426 1010
rect 3799 870 5150 970
rect 5250 870 5256 970
rect 3658 713 3664 722
rect 3653 679 3664 713
rect 3658 670 3664 679
rect 3716 670 3722 722
rect 3799 720 3899 870
rect 4326 840 4426 870
rect 4320 740 4326 840
rect 4426 740 4432 840
rect 4350 738 4402 740
rect 3824 719 3876 720
rect 3824 670 3876 673
rect 3978 670 3984 722
rect 4036 713 4042 722
rect 4036 679 4047 713
rect 4036 670 4042 679
rect 3800 630 3900 670
rect 4730 630 4829 636
rect 3800 530 4350 630
rect 4399 584 4730 630
rect 4400 531 4730 584
rect 4400 530 4829 531
rect 3658 293 3664 302
rect 3653 259 3664 293
rect 3658 250 3664 259
rect 3716 250 3722 302
rect 3800 300 3900 530
rect 4730 525 4829 530
rect 4350 476 4402 482
rect 4350 418 4402 424
rect 4359 413 4393 418
rect 3824 299 3876 300
rect 3824 250 3876 253
rect 3978 250 3984 302
rect 4036 293 4042 302
rect 4036 259 4047 293
rect 4036 250 4042 259
rect 3800 160 3900 250
rect 3794 60 3800 160
rect 3900 60 3906 160
rect 4320 -100 4420 -94
rect 3280 -190 3750 -100
rect 3500 -540 3750 -190
rect 3830 -540 4080 -100
rect 4170 -200 4320 -100
rect 4170 -540 4420 -200
rect 2120 -1770 2370 -1330
rect 2450 -1770 2700 -1330
rect 2780 -1770 3030 -1330
rect 3110 -1770 3360 -1330
rect 3670 -1770 3920 -1330
rect 4000 -1770 4250 -1330
<< via1 >>
rect 2770 2824 2870 2830
rect 2770 2736 2776 2824
rect 2776 2736 2864 2824
rect 2864 2736 2870 2824
rect 2770 2730 2870 2736
rect 4321 1980 4420 2079
rect 2100 870 2200 970
rect 3799 1720 3900 1820
rect 3659 1560 3711 1612
rect 3987 1560 4039 1612
rect 4210 1704 4310 1710
rect 4210 1616 4216 1704
rect 4216 1616 4304 1704
rect 4304 1616 4310 1704
rect 4210 1610 4310 1616
rect 4350 1377 4402 1429
rect 4530 1210 4630 1310
rect 3659 1120 3711 1172
rect 3987 1120 4039 1172
rect 4326 1010 4426 1110
rect 5150 870 5250 970
rect 3664 670 3716 722
rect 4326 740 4426 840
rect 3984 670 4036 722
rect 4730 531 4829 630
rect 3664 250 3716 302
rect 4350 424 4402 476
rect 3984 250 4036 302
rect 3800 60 3900 160
rect 4320 -200 4420 -100
<< metal2 >>
rect 4480 16620 4680 16820
rect 3160 16610 3260 16619
rect 4480 16610 4630 16620
rect 3260 16510 4630 16610
rect 3160 16501 3260 16510
rect 4530 2830 4630 16510
rect 2764 2730 2770 2830
rect 2870 2730 4630 2830
rect 4530 2079 4630 2730
rect 4315 1980 4321 2079
rect 4420 1980 4630 2079
rect 4530 1820 4630 1980
rect 3790 1720 3799 1820
rect 3900 1720 4630 1820
rect 4210 1710 4310 1720
rect 3530 1612 4060 1636
rect 3530 1560 3659 1612
rect 3711 1560 3987 1612
rect 4039 1560 4060 1612
rect 4210 1604 4310 1610
rect 3530 1536 4060 1560
rect 4530 1560 4630 1720
rect 3530 1196 3630 1536
rect 4530 1460 4829 1560
rect 4326 1429 4426 1460
rect 4326 1377 4350 1429
rect 4402 1377 4426 1429
rect 3530 1172 4060 1196
rect 3530 1120 3659 1172
rect 3711 1120 3987 1172
rect 4039 1120 4060 1172
rect 3530 1096 4060 1120
rect 4326 1110 4426 1377
rect 1390 970 1590 1020
rect 3530 970 3630 1096
rect 4326 1004 4426 1010
rect 4530 1310 4630 1316
rect 1390 870 2100 970
rect 2200 870 3630 970
rect 1390 820 1590 870
rect 3530 746 3630 870
rect 4326 840 4426 846
rect 3530 722 4060 746
rect 3530 670 3664 722
rect 3716 670 3984 722
rect 4036 670 4060 722
rect 3530 646 4060 670
rect 3530 326 3630 646
rect 4326 476 4426 740
rect 4326 424 4350 476
rect 4402 424 4426 476
rect 4326 400 4426 424
rect 3530 302 4060 326
rect 3530 250 3664 302
rect 3716 250 3984 302
rect 4036 250 4060 302
rect 3530 226 4060 250
rect 3800 160 3900 166
rect 4530 160 4630 1210
rect 4730 630 4829 1460
rect 5150 970 5350 1020
rect 5250 870 5350 970
rect 5150 820 5350 870
rect 4724 531 4730 630
rect 4829 531 4835 630
rect 3900 60 4630 160
rect 3800 54 3900 60
rect 4530 -100 4630 60
rect 4314 -200 4320 -100
rect 4420 -200 4630 -100
rect 4530 -3590 4630 -200
rect 4940 -3590 5040 -3581
rect 4530 -3690 4940 -3590
rect 4530 -3790 4630 -3690
rect 4940 -3699 5040 -3690
rect 4480 -3990 4680 -3790
<< via2 >>
rect 3160 16510 3260 16610
rect 4940 -3690 5040 -3590
<< metal3 >>
rect 3155 16610 3265 16615
rect 3155 16605 3160 16610
rect 3260 16605 3265 16610
rect 3155 16499 3265 16505
rect 4935 -3585 5045 -3579
rect 4935 -3690 4940 -3685
rect 5040 -3690 5045 -3685
rect 4935 -3695 5045 -3690
<< via3 >>
rect 3155 16510 3160 16605
rect 3160 16510 3260 16605
rect 3260 16510 3265 16605
rect 3155 16505 3265 16510
rect 4935 -3590 5045 -3585
rect 4935 -3685 4940 -3590
rect 4940 -3685 5040 -3590
rect 5040 -3685 5045 -3590
<< metal4 >>
rect 3150 16605 3270 16615
rect 3150 16505 3155 16605
rect 3265 16505 3270 16605
rect 3150 -3540 3270 16505
rect 4930 -3585 5050 16380
rect 4930 -3685 4935 -3585
rect 5045 -3685 5050 -3585
rect 4930 -3695 5050 -3685
use sky130_fd_pr__res_xhigh_po_0p35_UPT64K  sky130_fd_pr__res_xhigh_po_0p35_UPT64K_0 paramcells
timestamp 1718125978
transform 1 0 3960 0 1 2802
box -450 -982 450 982
use sky130_fd_pr__res_xhigh_po_0p35_UPT64K  sky130_fd_pr__res_xhigh_po_0p35_UPT64K_1
timestamp 1718125978
transform 1 0 3960 0 1 -948
box -450 -982 450 982
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC4 paramcells
timestamp 1713813547
transform 1 0 3346 0 1 6420
box -1686 -9960 1686 9960
use sky130_fd_pr__pfet_01v8_6QYSWZ  XM3 paramcells
timestamp 1713241921
transform 0 1 3849 -1 0 1146
box -226 -319 226 319
use sky130_fd_pr__nfet_01v8_723X3M  XM4 paramcells
timestamp 1712827999
transform 0 1 3850 -1 0 696
box -216 -310 216 310
use sky130_fd_pr__pfet_01v8_6QYSWZ  XM5
timestamp 1713241921
transform 0 1 3849 -1 0 1586
box -226 -319 226 319
use sky130_fd_pr__nfet_01v8_723X3M  XM6
timestamp 1712827999
transform 0 1 3850 -1 0 276
box -216 -310 216 310
use sky130_fd_pr__pfet_01v8_6QYSWZ  XM7
timestamp 1713241921
transform 1 0 4376 0 1 1239
box -226 -319 226 319
use sky130_fd_pr__nfet_01v8_723X3M  XM8
timestamp 1712827999
transform 1 0 4376 0 1 610
box -216 -310 216 310
use sky130_fd_pr__res_xhigh_po_0p35_J44QPS  XR3 paramcells
timestamp 1718125978
transform 1 0 2742 0 1 252
box -782 -2182 782 2182
<< labels >>
flabel metal2 1390 820 1590 1020 0 FreeSans 256 0 0 0 AIN
port 2 nsew
flabel metal2 5150 820 5350 1020 0 FreeSans 256 0 0 0 DOUT
port 3 nsew
flabel metal2 4480 16620 4680 16820 0 FreeSans 256 0 0 0 SG_DVDD
port 1 nsew
flabel metal2 4480 -3990 4680 -3790 0 FreeSans 256 0 0 0 SG_DVSS
port 4 nsew
flabel mvpsubdiff 4208 4445 4208 4445 0 FreeSans 320 0 0 0 VSUB
port 5 nsew
<< end >>
