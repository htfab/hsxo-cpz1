magic
tech sky130A
magscale 1 2
timestamp 1713812475
<< dnwell >>
rect -1970 -7210 5210 4580
rect -2520 -14610 2220 -9310
<< nwell >>
rect -2080 3960 5320 4690
rect -2080 3500 130 3960
rect -2080 -6990 -1764 3500
rect 5000 2760 5320 3960
rect 5004 -6890 5320 2760
rect 5000 -6990 5320 -6890
rect -2080 -7320 5320 -6990
rect -2600 -9782 2300 -9230
rect -2600 -12460 -1840 -9782
rect -2600 -14404 -2314 -12460
rect 1414 -14404 2300 -9782
rect -2600 -14690 2300 -14404
<< nsubdiff >>
rect -2563 -9287 2263 -9267
rect -2563 -9321 -2483 -9287
rect 2183 -9321 2263 -9287
rect -2563 -9341 2263 -9321
rect -2563 -9347 -2489 -9341
rect -2563 -14573 -2543 -9347
rect -2509 -14573 -2489 -9347
rect -2563 -14579 -2489 -14573
rect 2189 -9347 2263 -9341
rect 2189 -14573 2209 -9347
rect 2243 -14573 2263 -9347
rect 2189 -14579 2263 -14573
rect -2563 -14599 2263 -14579
rect -2563 -14633 -2483 -14599
rect 2183 -14633 2263 -14599
rect -2563 -14653 2263 -14633
<< mvnsubdiff >>
rect -2013 4603 5253 4623
rect -2013 4569 -1933 4603
rect 5173 4569 5253 4603
rect -2013 4549 5253 4569
rect -2013 4543 -1939 4549
rect -2013 -7173 -1993 4543
rect -1959 -7173 -1939 4543
rect -2013 -7179 -1939 -7173
rect 5179 4543 5253 4549
rect 5179 -7173 5199 4543
rect 5233 -7173 5253 4543
rect 5179 -7179 5253 -7173
rect -2013 -7199 5253 -7179
rect -2013 -7233 -1933 -7199
rect 5173 -7233 5253 -7199
rect -2013 -7253 5253 -7233
<< nsubdiffcont >>
rect -2483 -9321 2183 -9287
rect -2543 -14573 -2509 -9347
rect 2209 -14573 2243 -9347
rect -2483 -14633 2183 -14599
<< mvnsubdiffcont >>
rect -1933 4569 5173 4603
rect -1993 -7173 -1959 4543
rect 5199 -7173 5233 4543
rect -1933 -7233 5173 -7199
<< locali >>
rect -1993 4569 -1933 4603
rect 5173 4569 5233 4603
rect -1993 4543 -1959 4569
rect -1993 -7199 -1959 -7173
rect 5199 4543 5233 4569
rect 5199 -7199 5233 -7173
rect -1993 -7233 -1933 -7199
rect 5173 -7233 5233 -7199
rect -2543 -9321 -2483 -9287
rect 2183 -9321 2243 -9287
rect -2543 -9347 -2509 -9321
rect -2543 -14599 -2509 -14573
rect 2209 -9347 2243 -9321
rect 2209 -14599 2243 -14573
rect -2543 -14633 -2483 -14599
rect 2183 -14633 2243 -14599
rect 4587 -14963 4993 -14557
<< metal1 >>
rect 2520 6340 3320 6346
rect 3320 5540 5794 6340
rect 2520 5534 3320 5540
rect 540 4630 740 4830
rect 4994 3632 5794 5540
rect -3940 -8960 -3740 -7560
rect -3510 -8960 -3310 -7570
rect -3090 -8570 -2890 -7560
rect -2670 -8570 -2470 -7560
rect -2270 -7770 -2070 -7570
rect -1850 -7760 -1650 -7560
rect 1246 -8570 1446 -8564
rect -3096 -8770 -3090 -8570
rect -2890 -8770 -2884 -8570
rect -2670 -8770 1246 -8570
rect 1246 -8776 1446 -8770
rect -3946 -9160 -3940 -8960
rect -3740 -9160 -3734 -8960
rect -3510 -9160 -1014 -8960
rect -814 -9160 -808 -8960
rect -3409 -11803 -3403 -11397
rect -2997 -11803 -2991 -11397
rect -3403 -14767 -2997 -11803
rect 4587 -14557 4993 -14551
rect -3403 -14963 4587 -14767
rect -3403 -15173 4993 -14963
<< via1 >>
rect 2520 5540 3320 6340
rect -3090 -8770 -2890 -8570
rect 1246 -8770 1446 -8570
rect -3940 -9160 -3740 -8960
rect -1014 -9160 -814 -8960
rect -3403 -11803 -2997 -11397
rect 4587 -14963 4993 -14557
<< metal2 >>
rect 2520 6340 3320 6349
rect -3946 5540 780 6340
rect 1580 5540 1589 6340
rect 2514 5540 2520 6340
rect 3320 5540 3326 6340
rect -3946 4430 -3146 5540
rect 2520 5531 3320 5540
rect -3950 3630 -3146 4430
rect -3946 3626 -3146 3630
rect 2694 3626 3494 4430
rect 5800 -2300 6600 -1500
rect 5800 -3560 6600 -2760
rect 5800 -4840 6600 -4040
rect 5800 -6130 6600 -5330
rect -3146 -6560 -2346 -6555
rect -3150 -7360 -2346 -6560
rect -3146 -7373 -2346 -7360
rect -3090 -8570 -2890 -8564
rect -2890 -8770 -274 -8570
rect 1240 -8770 1246 -8570
rect 1446 -8770 1452 -8570
rect -3090 -8776 -2890 -8770
rect -3940 -8960 -3740 -8954
rect -1014 -8960 -814 -8954
rect -3740 -9160 -1754 -8960
rect -3940 -9166 -3740 -9160
rect -1954 -9530 -1754 -9160
rect -1014 -9536 -814 -9160
rect -474 -9530 -274 -8770
rect 1246 -9536 1446 -8770
rect -3403 -11397 -2997 -11391
rect -2920 -11397 -1954 -11394
rect -2997 -11800 -1954 -11397
rect -2997 -11803 -2427 -11800
rect -3403 -11809 -2997 -11803
rect -2360 -11806 -1960 -11800
rect 2300 -12480 2700 -12080
rect 2300 -13070 2700 -12670
rect 2500 -13490 2700 -13290
rect -2560 -14170 -1960 -13770
rect 3690 -14110 6760 -13710
rect -2560 -14770 -2160 -14170
rect 3690 -14770 4090 -14110
rect 4587 -14551 4993 -14548
rect 6360 -14550 6760 -14110
rect -2560 -15170 4090 -14770
rect 4575 -14557 5005 -14551
rect 4575 -14957 4587 -14557
rect 4581 -14963 4587 -14957
rect 4993 -14957 5005 -14557
rect 4993 -14963 4999 -14957
rect 6360 -14959 6760 -14950
rect 4587 -14972 4993 -14963
<< via2 >>
rect 780 5540 1580 6340
rect 2520 5540 3320 6340
rect 4587 -14963 4993 -14557
rect 6360 -14950 6760 -14550
<< metal3 >>
rect 755 6355 1575 6365
rect 755 5555 765 6355
rect 2515 6345 3325 6355
rect 1575 6340 1585 6345
rect 765 5549 780 5555
rect 775 5540 780 5549
rect 1580 5540 1585 6340
rect 775 5535 1070 5540
rect 1065 5475 1070 5535
rect 1275 5535 1585 5540
rect 2515 5529 2831 5535
rect 2825 5481 2831 5529
rect 3029 5529 3325 5535
rect 3029 5481 3035 5529
rect 2830 5480 3030 5481
rect 1065 5469 1275 5475
rect 6355 -14540 6765 -14539
rect 6342 -14545 6765 -14540
rect 6342 -14546 6355 -14545
rect 4582 -14552 4998 -14546
rect 4575 -14565 4582 -14559
rect 4993 -14963 4998 -14958
rect 6760 -14950 6765 -14945
rect 6758 -14952 6765 -14950
rect 6342 -14955 6765 -14952
rect 6342 -14962 6758 -14955
rect 4985 -14965 4998 -14963
rect 4575 -14968 4998 -14965
rect 4575 -14975 4985 -14968
<< via3 >>
rect 765 6340 1575 6355
rect 765 5555 780 6340
rect 780 5555 1575 6340
rect 1070 5540 1275 5555
rect 1070 5475 1275 5540
rect 2515 6340 3325 6345
rect 2515 5540 2520 6340
rect 2520 5540 3320 6340
rect 3320 5540 3325 6340
rect 2515 5535 3325 5540
rect 2831 5481 3029 5535
rect 6355 -14546 6765 -14545
rect 4582 -14557 4998 -14552
rect 4582 -14565 4587 -14557
rect 4575 -14963 4587 -14565
rect 4587 -14958 4993 -14557
rect 4993 -14958 4998 -14557
rect 4587 -14963 4985 -14958
rect 6342 -14550 6765 -14546
rect 6342 -14950 6360 -14550
rect 6360 -14945 6760 -14550
rect 6760 -14945 6765 -14550
rect 6360 -14950 6758 -14945
rect 6342 -14952 6758 -14950
rect 4575 -14965 4985 -14963
<< metal4 >>
rect 764 6355 1576 6356
rect 764 5555 765 6355
rect 1575 5555 1576 6355
rect 764 5554 1070 5555
rect 1060 5475 1070 5554
rect 1275 5554 1576 5555
rect 2514 6345 3326 6346
rect 1275 5475 1280 5554
rect 2514 5535 2515 6345
rect 3325 5535 3326 6345
rect 2514 5534 2831 5535
rect 1060 5470 1280 5475
rect 2830 5481 2831 5534
rect 3029 5534 3326 5535
rect 3029 5481 3030 5534
rect 1070 -14530 1270 5470
rect 2830 -14540 3030 5481
rect 4675 -14551 4875 5410
rect 6450 -14544 6650 5410
rect 6354 -14545 6766 -14544
rect 6341 -14546 6355 -14545
rect 4581 -14552 4999 -14551
rect 4581 -14564 4582 -14552
rect 4574 -14565 4582 -14564
rect 4574 -14965 4575 -14565
rect 4998 -14958 4999 -14552
rect 6341 -14952 6342 -14546
rect 6765 -14945 6766 -14545
rect 6758 -14946 6766 -14945
rect 6758 -14952 6759 -14946
rect 6341 -14953 6759 -14952
rect 4985 -14959 4999 -14958
rect 4985 -14965 4986 -14959
rect 4574 -14966 4986 -14965
rect 4579 -14971 4981 -14966
use power_gating_ad  power_gating_ad_1
timestamp 1713809040
transform 1 0 -2356 0 1 896
box -1594 -8666 8950 3936
use power_gating_dd  power_gating_dd_0
timestamp 1713804741
transform 1 0 -3664 0 1 -8010
box 1304 -6360 6360 -1320
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC3
timestamp 1713804741
transform 1 0 1296 0 1 -4550
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC4
timestamp 1713804741
transform 1 0 4916 0 1 -4550
box -1686 -9960 1686 9960
<< labels >>
flabel metal2 -3940 -9160 -3740 -8960 0 FreeSans 256 0 0 0 ENA
port 9 nsew
flabel via1 -3090 -8770 -2890 -8570 0 FreeSans 256 0 0 0 STDBY
port 12 nsew
flabel metal2 -2360 -11800 -1960 -11400 0 FreeSans 256 0 0 0 DVDD
port 3 nsew
flabel metal2 2300 -13070 2700 -12670 0 FreeSans 256 0 0 0 SG_DVSS
port 10 nsew
flabel metal2 2300 -12480 2700 -12080 0 FreeSans 256 0 0 0 SG_DVDD
port 5 nsew
flabel metal2 -3950 3630 -3150 4430 0 FreeSans 256 0 0 0 AVDD
port 6 nsew
flabel metal1 -1850 -7760 -1650 -7560 0 FreeSans 256 0 0 0 XIN
port 16 nsew
flabel metal1 -2270 -7770 -2070 -7570 0 FreeSans 256 0 0 0 EG_IBIAS
port 4 nsew
flabel metal1 540 4630 740 4830 0 FreeSans 256 0 0 0 IBIAS
port 7 nsew
flabel metal2 5800 -3560 6600 -2760 0 FreeSans 256 0 0 0 EG_AVDD
port 8 nsew
flabel metal2 5800 -4840 6600 -4040 0 FreeSans 256 0 0 0 EG_AVSS
port 13 nsew
flabel metal2 5800 -6130 6600 -5330 0 FreeSans 256 0 0 0 SG_AVSS
port 11 nsew
flabel metal2 5800 -2300 6600 -1500 0 FreeSans 256 0 0 0 SG_AVDD
port 2 nsew
flabel metal2 2500 -13490 2700 -13290 0 FreeSans 256 0 0 0 DOUT
port 1 nsew
flabel metal2 -2360 -14170 -1960 -13770 0 FreeSans 256 0 0 0 DVSS
port 15 nsew
flabel metal2 -3150 -7360 -2350 -6560 0 FreeSans 256 0 0 0 AVSS
port 14 nsew
<< end >>
