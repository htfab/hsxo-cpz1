magic
tech sky130A
magscale 1 2
timestamp 1718126023
<< dnwell >>
rect 380 330 9870 15250
rect 11130 4760 13440 15250
<< nwell >>
rect 270 14640 9980 15360
rect 270 12480 1500 14640
rect 270 536 586 12480
rect 9050 7650 9980 14640
rect 9664 536 9980 7650
rect 11020 6470 13550 15360
rect 11020 4966 11336 6470
rect 13234 4966 13550 6470
rect 11020 4650 13550 4966
rect 270 220 9980 536
<< mvpsubdiff >>
rect 9030 3990 9430 4014
rect 9030 2966 9430 2990
rect 12650 6180 13050 6204
rect 12650 5156 13050 5180
<< mvnsubdiff >>
rect 337 15273 9913 15293
rect 337 15239 417 15273
rect 9833 15239 9913 15273
rect 337 15219 9913 15239
rect 337 15213 411 15219
rect 337 367 357 15213
rect 391 367 411 15213
rect 9839 15213 9913 15219
rect 1070 13570 1470 13594
rect 1070 12546 1470 12570
rect 337 361 411 367
rect 9839 367 9859 15213
rect 9893 367 9913 15213
rect 11087 15273 13483 15293
rect 11087 15239 11167 15273
rect 13403 15239 13483 15273
rect 11087 15219 13483 15239
rect 11087 15213 11161 15219
rect 11087 4797 11107 15213
rect 11141 4797 11161 15213
rect 13409 15213 13483 15219
rect 12050 7560 12450 7584
rect 12050 6536 12450 6560
rect 11087 4791 11161 4797
rect 13409 4797 13429 15213
rect 13463 4797 13483 15213
rect 13409 4791 13483 4797
rect 11087 4771 13483 4791
rect 11087 4737 11167 4771
rect 13403 4737 13483 4771
rect 11087 4717 13483 4737
rect 9839 361 9913 367
rect 337 341 9913 361
rect 337 307 417 341
rect 9833 307 9913 341
rect 337 287 9913 307
<< mvpsubdiffcont >>
rect 9030 2990 9430 3990
rect 12650 5180 13050 6180
<< mvnsubdiffcont >>
rect 417 15239 9833 15273
rect 357 367 391 15213
rect 1070 12570 1470 13570
rect 9859 367 9893 15213
rect 11167 15239 13403 15273
rect 11107 4797 11141 15213
rect 12050 6560 12450 7560
rect 13429 4797 13463 15213
rect 11167 4737 13403 4771
rect 417 307 9833 341
<< locali >>
rect 357 15239 417 15273
rect 9833 15239 9893 15273
rect 357 15213 391 15239
rect 9859 15213 9893 15239
rect 1518 14472 9032 14626
rect 1070 13570 1470 13586
rect 1518 13570 1672 14472
rect 1470 12570 1672 13570
rect 1070 12554 1470 12570
rect 976 12104 1130 12108
rect 1296 12104 1450 12108
rect 972 11950 1454 12104
rect 976 9590 1130 11950
rect 1296 9590 1450 11950
rect 976 9270 1450 9590
rect 976 7608 1130 9270
rect 1296 7608 1450 9270
rect 1518 7822 1672 12570
rect 6842 7822 7112 14472
rect 7858 7822 8132 14472
rect 8878 7822 9032 14472
rect 1518 7668 9032 7822
rect 938 7454 8992 7608
rect 938 822 1092 7454
rect 1364 822 1632 7454
rect 2378 822 2652 7454
rect 7822 822 8092 7454
rect 8838 3990 8992 7454
rect 9030 3990 9430 4006
rect 8838 2990 9030 3990
rect 8838 2808 8992 2990
rect 9030 2974 9430 2990
rect 8838 2768 9498 2808
rect 8838 2654 9538 2768
rect 8838 822 9112 2654
rect 9384 822 9538 2654
rect 938 708 9538 822
rect 938 668 9498 708
rect 357 341 391 367
rect 11107 15239 11167 15273
rect 13403 15239 13463 15273
rect 11107 15213 11141 15239
rect 13429 15213 13463 15239
rect 11758 14472 12812 14626
rect 11758 7822 11912 14472
rect 12658 7822 12812 14472
rect 11758 7668 12812 7822
rect 12050 7560 12450 7668
rect 12050 6544 12450 6560
rect 11718 6274 12298 6428
rect 11718 5242 11872 6274
rect 12144 6180 12298 6274
rect 12650 6180 13050 6196
rect 12144 5242 12650 6180
rect 11718 5180 12650 5242
rect 11718 5088 12298 5180
rect 12650 5164 13050 5180
rect 11107 4771 11141 4797
rect 13429 4771 13463 4797
rect 11107 4737 11167 4771
rect 13403 4737 13463 4771
rect 9859 341 9893 367
rect 357 307 417 341
rect 9833 307 9893 341
<< viali >>
rect 1070 12570 1470 13570
rect 9030 2990 9430 3990
rect 12050 6560 12450 7560
rect 12660 5210 13040 6150
<< metal1 >>
rect 1750 14380 9280 14580
rect 9480 14380 12590 14580
rect 1058 13570 1482 13576
rect 1058 12570 1070 13570
rect 1470 12570 1482 13570
rect 1058 12564 1482 12570
rect 1665 12140 1671 12940
rect 1787 12140 1793 12940
rect 1981 12140 1987 12940
rect 2103 12140 2109 12940
rect 2297 12140 2303 12940
rect 2419 12140 2425 12940
rect 2613 12140 2619 12940
rect 2735 12140 2741 12940
rect 2929 12140 2935 12940
rect 3051 12140 3057 12940
rect 3245 12140 3251 12940
rect 3367 12140 3373 12940
rect 3561 12140 3567 12940
rect 3683 12140 3689 12940
rect 3877 12140 3883 12940
rect 3999 12140 4005 12940
rect 4193 12140 4199 12940
rect 4315 12140 4321 12940
rect 4509 12140 4515 12940
rect 4631 12140 4637 12940
rect 4825 12140 4831 12940
rect 4947 12140 4953 12940
rect 5141 12140 5147 12940
rect 5263 12140 5269 12940
rect 5457 12140 5463 12940
rect 5579 12140 5585 12940
rect 5773 12140 5779 12940
rect 5895 12140 5901 12940
rect 6089 12140 6095 12940
rect 6211 12140 6217 12940
rect 6405 12140 6411 12940
rect 6527 12140 6533 12940
rect 6721 12140 6727 12940
rect 6843 12140 6849 12940
rect 7105 12140 7111 12940
rect 7227 12140 7233 12940
rect 7421 12140 7427 12940
rect 7543 12140 7549 12940
rect 7737 12140 7743 12940
rect 7859 12140 7865 12940
rect 8125 12140 8131 12940
rect 8247 12140 8253 12940
rect 8441 12140 8447 12940
rect 8563 12140 8569 12940
rect 8757 12140 8763 12940
rect 8879 12140 8885 12940
rect 11905 12140 11911 12940
rect 12027 12140 12033 12940
rect 12221 12140 12227 12940
rect 12343 12140 12349 12940
rect 12537 12140 12543 12940
rect 12659 12140 12665 12940
rect 1113 11910 1313 11916
rect 1113 11454 1313 11460
rect 1113 9830 1313 10080
rect 1823 9950 1829 10150
rect 1945 9950 1951 10150
rect 2139 9950 2145 10150
rect 2261 9950 2267 10150
rect 2455 9950 2461 10150
rect 2577 9950 2583 10150
rect 2771 9950 2777 10150
rect 2893 9950 2899 10150
rect 3087 9950 3093 10150
rect 3209 9950 3215 10150
rect 3403 9950 3409 10150
rect 3525 9950 3531 10150
rect 3719 9950 3725 10150
rect 3841 9950 3847 10150
rect 4035 9950 4041 10150
rect 4157 9950 4163 10150
rect 4351 9950 4357 10150
rect 4473 9950 4479 10150
rect 4667 9950 4673 10150
rect 4789 9950 4795 10150
rect 4983 9950 4989 10150
rect 5105 9950 5111 10150
rect 5299 9950 5305 10150
rect 5421 9950 5427 10150
rect 5615 9950 5621 10150
rect 5737 9950 5743 10150
rect 5931 9950 5937 10150
rect 6053 9950 6059 10150
rect 6247 9950 6253 10150
rect 6369 9950 6375 10150
rect 6563 9950 6569 10150
rect 6685 9950 6691 10150
rect 7263 9950 7269 10150
rect 7385 9950 7391 10150
rect 7579 9950 7585 10150
rect 7701 9950 7707 10150
rect 8283 9950 8289 10150
rect 8405 9950 8411 10150
rect 8599 9950 8605 10150
rect 8721 9950 8727 10150
rect 12063 9950 12069 10150
rect 12185 9950 12191 10150
rect 12379 9950 12385 10150
rect 12501 9950 12507 10150
rect 680 9630 1313 9830
rect 680 7940 880 9630
rect 1113 9230 1313 9236
rect 1113 8784 1313 8790
rect 360 7740 880 7940
rect -30 4300 170 4306
rect -30 110 170 4100
rect 360 3150 560 7740
rect 1113 7570 1313 8230
rect 1740 7710 7650 7910
rect 7850 7710 12590 7910
rect 724 7370 730 7570
rect 930 7370 1313 7570
rect 1700 7370 7750 7570
rect 8160 7370 9770 7570
rect 12038 7560 12462 7566
rect 12038 7430 12050 7560
rect 360 480 560 2950
rect 730 910 930 7370
rect 1085 5130 1091 5330
rect 1207 5130 1213 5330
rect 1625 5130 1631 5330
rect 1747 5130 1753 5330
rect 1941 5130 1947 5330
rect 2063 5130 2069 5330
rect 2257 5130 2263 5330
rect 2379 5130 2385 5330
rect 2645 5130 2651 5330
rect 2767 5130 2773 5330
rect 2961 5130 2967 5330
rect 3083 5130 3089 5330
rect 3277 5130 3283 5330
rect 3399 5130 3405 5330
rect 3593 5130 3599 5330
rect 3715 5130 3721 5330
rect 3909 5130 3915 5330
rect 4031 5130 4037 5330
rect 4225 5130 4231 5330
rect 4347 5130 4353 5330
rect 4541 5130 4547 5330
rect 4663 5130 4669 5330
rect 4857 5130 4863 5330
rect 4979 5130 4985 5330
rect 5173 5130 5179 5330
rect 5295 5130 5301 5330
rect 5489 5130 5495 5330
rect 5611 5130 5617 5330
rect 5805 5130 5811 5330
rect 5927 5130 5933 5330
rect 6121 5130 6127 5330
rect 6243 5130 6249 5330
rect 6437 5130 6443 5330
rect 6559 5130 6565 5330
rect 6753 5130 6759 5330
rect 6875 5130 6881 5330
rect 7069 5130 7075 5330
rect 7191 5130 7197 5330
rect 7385 5130 7391 5330
rect 7507 5130 7513 5330
rect 7701 5130 7707 5330
rect 7823 5130 7829 5330
rect 8085 5130 8091 5330
rect 8207 5130 8213 5330
rect 8401 5130 8407 5330
rect 8523 5130 8529 5330
rect 8717 5130 8723 5330
rect 8839 5130 8845 5330
rect 9018 3990 9442 3996
rect 1243 2950 1249 3750
rect 1365 2950 1371 3750
rect 1783 2950 1789 3750
rect 1905 2950 1911 3750
rect 2099 2950 2105 3750
rect 2221 2950 2227 3750
rect 2803 2950 2809 3150
rect 2925 2950 2931 3150
rect 3119 2950 3125 3150
rect 3241 2950 3247 3150
rect 3435 2950 3441 3150
rect 3557 2950 3563 3150
rect 3751 2950 3757 3150
rect 3873 2950 3879 3150
rect 4067 2950 4073 3150
rect 4189 2950 4195 3150
rect 4383 2950 4389 3150
rect 4505 2950 4511 3150
rect 4699 2950 4705 3150
rect 4821 2950 4827 3150
rect 5015 2950 5021 3150
rect 5137 2950 5143 3150
rect 5331 2950 5337 3150
rect 5453 2950 5459 3150
rect 5647 2950 5653 3150
rect 5769 2950 5775 3150
rect 5963 2950 5969 3150
rect 6085 2950 6091 3150
rect 6279 2950 6285 3150
rect 6401 2950 6407 3150
rect 6595 2950 6601 3150
rect 6717 2950 6723 3150
rect 6911 2950 6917 3150
rect 7033 2950 7039 3150
rect 7227 2950 7233 3150
rect 7349 2950 7355 3150
rect 7543 2950 7549 3150
rect 7665 2950 7671 3150
rect 8243 2950 8249 3750
rect 8365 2950 8371 3750
rect 8559 2950 8565 3750
rect 8681 2950 8687 3750
rect 9018 2990 9030 3990
rect 9430 2990 9442 3990
rect 9018 2984 9442 2990
rect 9150 2770 9350 2780
rect 9570 2770 9770 7370
rect 10874 6630 10880 7430
rect 11680 6630 12050 7430
rect 12038 6560 12050 6630
rect 12450 6560 12462 7560
rect 12038 6554 12462 6560
rect 11460 6190 12080 6390
rect 11460 5330 11660 6190
rect 12650 6150 13050 6180
rect 11865 5866 11871 6066
rect 11987 5866 11993 6066
rect 12023 5410 12029 5770
rect 12145 5410 12151 5770
rect 11460 5130 12080 5330
rect 12650 5210 12660 6150
rect 13040 5210 13050 6150
rect 12650 5180 13050 5210
rect 11460 4960 11660 5130
rect 10754 4760 10760 4960
rect 10960 4760 11660 4960
rect 9144 2570 9150 2770
rect 9350 2570 9770 2770
rect 9570 2170 9770 2180
rect 9105 1970 9111 2170
rect 9227 1970 9233 2170
rect 9263 1310 9269 1510
rect 9385 1310 9391 1510
rect 9570 910 9770 1970
rect 730 710 1100 910
rect 1300 710 1306 910
rect 1700 710 7760 910
rect 8160 710 9770 910
rect 1700 480 1900 710
rect 360 280 1900 480
rect -30 -90 2230 110
rect 2030 -2196 2230 -90
rect 2030 -2402 2230 -2396
rect 3080 -2201 3280 710
rect 3080 -2407 3280 -2401
rect 4930 -2201 5130 710
rect 4930 -2407 5130 -2401
rect 9570 -3230 9770 710
rect 11180 -1740 13660 -1540
rect 13860 -1740 13866 -1540
rect 11180 -2190 11380 -1740
rect 11180 -2396 11380 -2390
<< via1 >>
rect 9280 14380 9480 14580
rect 1130 12730 1410 13420
rect 1671 12140 1787 12940
rect 1987 12140 2103 12940
rect 2303 12140 2419 12940
rect 2619 12140 2735 12940
rect 2935 12140 3051 12940
rect 3251 12140 3367 12940
rect 3567 12140 3683 12940
rect 3883 12140 3999 12940
rect 4199 12140 4315 12940
rect 4515 12140 4631 12940
rect 4831 12140 4947 12940
rect 5147 12140 5263 12940
rect 5463 12140 5579 12940
rect 5779 12140 5895 12940
rect 6095 12140 6211 12940
rect 6411 12140 6527 12940
rect 6727 12140 6843 12940
rect 7111 12140 7227 12940
rect 7427 12140 7543 12940
rect 7743 12140 7859 12940
rect 8131 12140 8247 12940
rect 8447 12140 8563 12940
rect 8763 12140 8879 12940
rect 11911 12140 12027 12940
rect 12227 12140 12343 12940
rect 12543 12140 12659 12940
rect 1113 11460 1313 11910
rect 1829 9950 1945 10150
rect 2145 9950 2261 10150
rect 2461 9950 2577 10150
rect 2777 9950 2893 10150
rect 3093 9950 3209 10150
rect 3409 9950 3525 10150
rect 3725 9950 3841 10150
rect 4041 9950 4157 10150
rect 4357 9950 4473 10150
rect 4673 9950 4789 10150
rect 4989 9950 5105 10150
rect 5305 9950 5421 10150
rect 5621 9950 5737 10150
rect 5937 9950 6053 10150
rect 6253 9950 6369 10150
rect 6569 9950 6685 10150
rect 7269 9950 7385 10150
rect 7585 9950 7701 10150
rect 8289 9950 8405 10150
rect 8605 9950 8721 10150
rect 12069 9950 12185 10150
rect 12385 9950 12501 10150
rect 1113 8790 1313 9230
rect -30 4100 170 4300
rect 7650 7710 7850 7910
rect 730 7370 930 7570
rect 360 2950 560 3150
rect 1091 5130 1207 5330
rect 1631 5130 1747 5330
rect 1947 5130 2063 5330
rect 2263 5130 2379 5330
rect 2651 5130 2767 5330
rect 2967 5130 3083 5330
rect 3283 5130 3399 5330
rect 3599 5130 3715 5330
rect 3915 5130 4031 5330
rect 4231 5130 4347 5330
rect 4547 5130 4663 5330
rect 4863 5130 4979 5330
rect 5179 5130 5295 5330
rect 5495 5130 5611 5330
rect 5811 5130 5927 5330
rect 6127 5130 6243 5330
rect 6443 5130 6559 5330
rect 6759 5130 6875 5330
rect 7075 5130 7191 5330
rect 7391 5130 7507 5330
rect 7707 5130 7823 5330
rect 8091 5130 8207 5330
rect 8407 5130 8523 5330
rect 8723 5130 8839 5330
rect 1249 2950 1365 3750
rect 1789 2950 1905 3750
rect 2105 2950 2221 3750
rect 2809 2950 2925 3150
rect 3125 2950 3241 3150
rect 3441 2950 3557 3150
rect 3757 2950 3873 3150
rect 4073 2950 4189 3150
rect 4389 2950 4505 3150
rect 4705 2950 4821 3150
rect 5021 2950 5137 3150
rect 5337 2950 5453 3150
rect 5653 2950 5769 3150
rect 5969 2950 6085 3150
rect 6285 2950 6401 3150
rect 6601 2950 6717 3150
rect 6917 2950 7033 3150
rect 7233 2950 7349 3150
rect 7549 2950 7665 3150
rect 8249 2950 8365 3750
rect 8565 2950 8681 3750
rect 9090 3150 9370 3850
rect 10880 6630 11680 7430
rect 11871 5866 11987 6066
rect 12029 5410 12145 5770
rect 12700 5300 13000 6060
rect 10760 4760 10960 4960
rect 9150 2570 9350 2770
rect 9111 1970 9227 2170
rect 9570 1970 9770 2170
rect 9269 1310 9385 1510
rect 1100 710 1300 910
rect 2030 -2396 2230 -2196
rect 3080 -2401 3280 -2201
rect 4930 -2401 5130 -2201
rect 13660 -1740 13860 -1540
rect 11180 -2390 11380 -2190
<< metal2 >>
rect 11880 18830 12680 18839
rect 8270 18810 9070 18819
rect 12680 18030 13570 18830
rect 11880 18021 12680 18030
rect 870 13420 1670 13570
rect 870 12940 1130 13420
rect -340 12730 1130 12940
rect 1410 12940 1670 13420
rect 8270 12940 9070 18010
rect 1410 12730 1671 12940
rect -340 12140 1671 12730
rect 1787 12140 1987 12940
rect 2103 12140 2303 12940
rect 2419 12140 2619 12940
rect 2735 12140 2935 12940
rect 3051 12140 3251 12940
rect 3367 12140 3567 12940
rect 3683 12140 3883 12940
rect 3999 12140 4199 12940
rect 4315 12140 4515 12940
rect 4631 12140 4831 12940
rect 4947 12140 5147 12940
rect 5263 12140 5463 12940
rect 5579 12140 5779 12940
rect 5895 12140 6095 12940
rect 6211 12140 6411 12940
rect 6527 12140 6727 12940
rect 6843 12140 7111 12940
rect 7227 12140 7427 12940
rect 7543 12140 7743 12940
rect 7859 12140 8131 12940
rect 8247 12140 8447 12940
rect 8563 12140 8763 12940
rect 8879 12140 9070 12940
rect 9280 14580 9480 14586
rect 1107 11460 1113 11910
rect 1313 11460 1319 11910
rect 1113 11260 1313 11460
rect 1113 11060 7280 11260
rect 7080 10150 7280 11060
rect 9280 10150 9480 14380
rect 12770 12940 13570 18030
rect 1630 9950 1829 10150
rect 1945 9950 2145 10150
rect 2261 9950 2461 10150
rect 2577 9950 2777 10150
rect 2893 9950 3093 10150
rect 3209 9950 3409 10150
rect 3525 9950 3725 10150
rect 3841 9950 4041 10150
rect 4157 9950 4357 10150
rect 4473 9950 4673 10150
rect 4789 9950 4989 10150
rect 5105 9950 5305 10150
rect 5421 9950 5621 10150
rect 5737 9950 5937 10150
rect 6053 9950 6253 10150
rect 6369 9950 6569 10150
rect 6685 9950 6870 10150
rect 7080 9950 7269 10150
rect 7385 9950 7585 10150
rect 7701 9950 7890 10150
rect 8100 9950 8289 10150
rect 8405 9950 8605 10150
rect 8721 9950 9480 10150
rect 10880 12140 11911 12940
rect 12027 12140 12227 12940
rect 12343 12140 12543 12940
rect 12659 12140 14360 12940
rect 1630 9230 1830 9950
rect 7080 9540 7280 9950
rect 8100 9540 8300 9950
rect 1107 8790 1113 9230
rect 1313 9030 1830 9230
rect 2210 9340 7280 9540
rect 7650 9340 8300 9540
rect 1313 8790 1319 9030
rect 730 7570 930 7576
rect -340 7370 730 7570
rect 730 7364 930 7370
rect 1113 5330 1313 8790
rect 2210 5330 2410 9340
rect 7650 7910 7850 9340
rect 7650 5330 7850 7710
rect 10880 7430 11680 12140
rect 11880 9950 12069 10150
rect 12185 9950 12385 10150
rect 12501 9950 12690 10150
rect 10880 6624 11680 6630
rect 12230 8460 12430 9950
rect 12230 8260 14356 8460
rect 12230 6066 12430 8260
rect 11620 5866 11871 6066
rect 11987 5866 12430 6066
rect 12640 6060 13440 6180
rect 12640 5770 12700 6060
rect 11070 5410 12029 5770
rect 12145 5410 12700 5770
rect -340 5130 1091 5330
rect 1207 5130 1400 5330
rect 1600 5130 1631 5330
rect 1747 5130 1947 5330
rect 2063 5130 2263 5330
rect 2379 5130 2410 5330
rect 2620 5130 2651 5330
rect 2767 5130 2967 5330
rect 3083 5130 3283 5330
rect 3399 5130 3599 5330
rect 3715 5130 3915 5330
rect 4031 5130 4231 5330
rect 4347 5130 4547 5330
rect 4663 5130 4863 5330
rect 4979 5130 5179 5330
rect 5295 5130 5495 5330
rect 5611 5130 5811 5330
rect 5927 5130 6127 5330
rect 6243 5130 6443 5330
rect 6559 5130 6759 5330
rect 6875 5130 7075 5330
rect 7191 5130 7391 5330
rect 7507 5130 7707 5330
rect 7823 5130 7850 5330
rect 8060 5130 8091 5330
rect 8207 5130 8407 5330
rect 8523 5130 8723 5330
rect 8839 5130 8870 5330
rect 12640 5300 12700 5410
rect 13000 5300 13440 6060
rect 1600 4300 1800 5130
rect -36 4100 -30 4300
rect 170 4100 1800 4300
rect 8060 4160 8260 5130
rect 7660 3960 8260 4160
rect 10760 4960 10960 4966
rect 40 2950 360 3150
rect 560 2950 566 3150
rect 1060 2950 1249 3750
rect 1365 2950 1789 3750
rect 1905 2950 2105 3750
rect 2221 2950 2410 3750
rect 7660 3150 7860 3960
rect 8830 3850 9630 3990
rect 8830 3750 9090 3850
rect 8070 3150 8249 3750
rect 2620 2950 2809 3150
rect 2925 2950 3125 3150
rect 3241 2950 3441 3150
rect 3557 2950 3757 3150
rect 3873 2950 4073 3150
rect 4189 2950 4389 3150
rect 4505 2950 4705 3150
rect 4821 2950 5021 3150
rect 5137 2950 5337 3150
rect 5453 2950 5653 3150
rect 5769 2950 5969 3150
rect 6085 2950 6285 3150
rect 6401 2950 6601 3150
rect 6717 2950 6917 3150
rect 7033 2950 7233 3150
rect 7349 2950 7549 3150
rect 7665 2950 7860 3150
rect 8060 2950 8249 3150
rect 8365 2950 8565 3750
rect 8681 3150 9090 3750
rect 9370 3150 9630 3850
rect 8681 2950 9630 3150
rect 1610 2110 2410 2950
rect 8070 2110 8870 2950
rect 9150 2770 9350 2776
rect 9150 2170 9350 2570
rect -340 1510 8870 2110
rect 9080 1970 9111 2170
rect 9227 1970 9570 2170
rect 9770 1970 10050 2170
rect -340 1310 9269 1510
rect 9385 1310 10540 1510
rect 1100 910 1300 916
rect 1100 -2192 1300 710
rect 1100 -2201 1500 -2192
rect 2030 -2196 2230 -2187
rect 1100 -2401 1300 -2201
rect 2024 -2396 2030 -2196
rect 2230 -2396 2236 -2196
rect 2400 -2201 2800 1310
rect 3080 -2201 3280 -2192
rect 4930 -2201 5130 -2192
rect 6710 -2201 6910 1310
rect 8070 710 10540 1310
rect 9740 -2201 10540 710
rect 1300 -3340 1500 -2401
rect 2030 -2405 2230 -2396
rect 3074 -2401 3080 -2201
rect 3280 -2401 3286 -2201
rect 4924 -2401 4930 -2201
rect 5130 -2401 5136 -2201
rect 6701 -2401 6710 -2201
rect 6910 -2401 6920 -2201
rect 3080 -2410 3280 -2401
rect 4930 -2410 5130 -2401
rect 2400 -2529 2800 -2520
rect 10540 -2421 10549 -2221
rect 9740 -3010 10540 -3001
rect 10760 -3340 10960 4760
rect 12640 -2190 13440 5300
rect 13660 -1540 13860 8260
rect 13660 -1746 13860 -1740
rect 11171 -2390 11180 -2190
rect 11380 -2390 11389 -2190
rect 13440 -2990 14370 -2190
rect 12640 -2999 13440 -2990
rect 1300 -3540 10960 -3340
<< via2 >>
rect 8270 18010 9070 18810
rect 11880 18030 12680 18830
rect 1300 -2401 1500 -2201
rect 2030 -2396 2230 -2196
rect 2400 -2520 2800 -2201
rect 3080 -2401 3280 -2201
rect 4930 -2401 5130 -2201
rect 6710 -2401 6910 -2201
rect 9740 -3001 10540 -2201
rect 11180 -2390 11380 -2190
rect 12640 -2990 13440 -2190
<< metal3 >>
rect 11875 18835 12685 18841
rect 8265 18810 9075 18815
rect 8265 18805 8270 18810
rect 9070 18805 9075 18810
rect 11875 18030 11880 18035
rect 12680 18030 12685 18035
rect 11875 18025 12175 18030
rect 12385 18025 12685 18030
rect 12175 18019 12385 18025
rect 8265 17999 9075 18005
rect 12635 -2185 13445 -2179
rect 11175 -2190 11185 -2185
rect 1295 -2196 1505 -2190
rect 1295 -2401 1300 -2396
rect 1500 -2401 1505 -2396
rect 1295 -2406 1505 -2401
rect 2025 -2196 2235 -2191
rect 2025 -2201 2030 -2196
rect 2230 -2201 2235 -2196
rect 2025 -2407 2235 -2401
rect 2395 -2196 2805 -2190
rect 3075 -2196 3285 -2190
rect 3075 -2401 3080 -2396
rect 3280 -2401 3285 -2396
rect 3075 -2406 3285 -2401
rect 4925 -2196 5135 -2190
rect 4925 -2401 4930 -2396
rect 5130 -2401 5135 -2396
rect 4925 -2406 5135 -2401
rect 6705 -2196 6915 -2190
rect 6705 -2401 6710 -2396
rect 6910 -2401 6915 -2396
rect 6705 -2406 6915 -2401
rect 9735 -2196 10545 -2190
rect 2395 -2531 2805 -2525
rect 11175 -2390 11180 -2190
rect 11175 -2395 11185 -2390
rect 11385 -2395 11391 -2185
rect 12635 -2990 12640 -2985
rect 13440 -2990 13445 -2985
rect 12635 -2995 13445 -2990
rect 9735 -3001 9740 -2996
rect 10540 -3001 10545 -2996
rect 9735 -3006 10545 -3001
<< via3 >>
rect 11875 18830 12685 18835
rect 8265 18010 8270 18805
rect 8270 18010 9070 18805
rect 9070 18010 9075 18805
rect 11875 18035 11880 18830
rect 11880 18035 12680 18830
rect 12680 18035 12685 18830
rect 12175 18030 12385 18035
rect 12175 18025 12385 18030
rect 8265 18005 9075 18010
rect 11185 -2190 11385 -2185
rect 1295 -2201 1505 -2196
rect 1295 -2396 1300 -2201
rect 1300 -2396 1500 -2201
rect 1500 -2396 1505 -2201
rect 2025 -2396 2030 -2201
rect 2030 -2396 2230 -2201
rect 2230 -2396 2235 -2201
rect 2025 -2401 2235 -2396
rect 2395 -2201 2805 -2196
rect 2395 -2520 2400 -2201
rect 2400 -2520 2800 -2201
rect 2800 -2520 2805 -2201
rect 3075 -2201 3285 -2196
rect 3075 -2396 3080 -2201
rect 3080 -2396 3280 -2201
rect 3280 -2396 3285 -2201
rect 4925 -2201 5135 -2196
rect 4925 -2396 4930 -2201
rect 4930 -2396 5130 -2201
rect 5130 -2396 5135 -2201
rect 6705 -2201 6915 -2196
rect 6705 -2396 6710 -2201
rect 6710 -2396 6910 -2201
rect 6910 -2396 6915 -2201
rect 9735 -2201 10545 -2196
rect 2395 -2525 2805 -2520
rect 9735 -2996 9740 -2201
rect 9740 -2996 10540 -2201
rect 10540 -2996 10545 -2201
rect 11185 -2390 11380 -2190
rect 11380 -2390 11385 -2190
rect 11185 -2395 11385 -2390
rect 12635 -2190 13445 -2185
rect 12635 -2985 12640 -2190
rect 12640 -2985 13440 -2190
rect 13440 -2985 13445 -2190
<< metal4 >>
rect 11874 18835 12686 18836
rect 8264 18805 9076 18806
rect 8264 18005 8265 18805
rect 9075 18005 9076 18805
rect 11874 18035 11875 18835
rect 12685 18035 12686 18835
rect 11874 18034 12175 18035
rect 12174 18025 12175 18034
rect 12385 18034 12686 18035
rect 12385 18025 12386 18034
rect 12174 18024 12386 18025
rect 8264 18004 9076 18005
rect 1300 -2195 1500 17850
rect 3079 -1831 3282 17851
rect 3080 -2195 3280 -1831
rect 4930 -2195 5130 17850
rect 6710 -2195 6910 17850
rect 8563 -2070 8763 18004
rect 10340 -2195 10540 17850
rect 12180 -2070 12380 18024
rect 11184 -2185 11386 -2184
rect 11184 -2190 11185 -2185
rect 1294 -2196 1506 -2195
rect 1294 -2396 1295 -2196
rect 1505 -2396 1506 -2196
rect 2394 -2196 2806 -2195
rect 1294 -2397 1506 -2396
rect 2024 -2201 2236 -2200
rect 2024 -2401 2025 -2201
rect 2235 -2401 2236 -2201
rect 2024 -2402 2236 -2401
rect 2030 -3010 2230 -2402
rect 2394 -2525 2395 -2196
rect 2805 -2525 2806 -2196
rect 3074 -2196 3286 -2195
rect 3074 -2396 3075 -2196
rect 3285 -2396 3286 -2196
rect 3074 -2397 3286 -2396
rect 4924 -2196 5136 -2195
rect 4924 -2396 4925 -2196
rect 5135 -2396 5136 -2196
rect 4924 -2397 5136 -2396
rect 6704 -2196 6916 -2195
rect 6704 -2396 6705 -2196
rect 6915 -2396 6916 -2196
rect 6704 -2397 6916 -2396
rect 9734 -2196 10546 -2195
rect 2394 -2526 2806 -2525
rect 2400 -3241 2800 -2526
rect 9734 -2996 9735 -2196
rect 10545 -2996 10546 -2196
rect 11180 -2395 11185 -2190
rect 11385 -2395 11386 -2185
rect 11180 -2396 11386 -2395
rect 12634 -2185 13446 -2184
rect 11180 -2400 11385 -2396
rect 11180 -2860 11380 -2400
rect 11660 -2775 11860 -2645
rect 12634 -2775 12635 -2185
rect 9734 -2997 10546 -2996
rect 11660 -2975 12635 -2775
rect 11660 -3105 11860 -2975
rect 12634 -2985 12635 -2975
rect 13445 -2190 13446 -2185
rect 13955 -2190 14155 17850
rect 13445 -2390 14155 -2190
rect 13445 -2985 13446 -2390
rect 12634 -2986 13446 -2985
use sky130_fd_pr__cap_mim_m3_1_VCTT89  XC1 paramcells
timestamp 1713748097
transform 1 0 2266 0 1 -3011
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC2 paramcells
timestamp 1713813547
transform 1 0 1546 0 1 7890
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC3
timestamp 1713813547
transform 1 0 8806 0 1 7890
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC4
timestamp 1713813547
transform 1 0 12426 0 1 7890
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  XC7
timestamp 1713813547
transform 1 0 5176 0 1 7890
box -1686 -9960 1686 9960
use sky130_fd_pr__cap_mim_m3_1_VCTT89  XC8
timestamp 1713748097
transform 1 0 11426 0 1 -2875
box -386 -240 386 240
use sky130_fd_pr__pfet_g5v0d10v5_AQSVLT  XM9 paramcells
timestamp 1713747467
transform 1 0 4257 0 1 11147
box -2757 -3497 2757 3497
use sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH  XM10 paramcells
timestamp 1713747467
transform 1 0 7485 0 1 11147
box -545 -3497 545 3497
use sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH  XM11
timestamp 1713747467
transform 1 0 8505 0 1 11147
box -545 -3497 545 3497
use sky130_fd_pr__nfet_g5v0d10v5_JULQJE  XM12 paramcells
timestamp 1713747467
transform 1 0 2005 0 1 4138
box -515 -3458 515 3458
use sky130_fd_pr__nfet_g5v0d10v5_KDBUUD  XM13 paramcells
timestamp 1713747467
transform 1 0 1228 0 1 4138
box -278 -3458 278 3458
use sky130_fd_pr__nfet_g5v0d10v5_844AHT  XM14 paramcells
timestamp 1713747467
transform 1 0 5237 0 1 4138
box -2727 -3458 2727 3458
use sky130_fd_pr__nfet_g5v0d10v5_JULQJE  XM15
timestamp 1713747467
transform 1 0 8465 0 1 4138
box -515 -3458 515 3458
use sky130_fd_pr__nfet_g5v0d10v5_YNEQJ5  XM16 paramcells
timestamp 1713747467
transform 1 0 9248 0 1 1738
box -278 -1058 278 1058
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  XM17 paramcells
timestamp 1713747467
transform 1 0 12008 0 1 5758
box -278 -658 278 658
use sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH  XM18
timestamp 1713747467
transform 1 0 12285 0 1 11147
box -545 -3497 545 3497
use sky130_fd_pr__res_xhigh_po_0p35_GPPFXN  XR1 paramcells
timestamp 1718126023
transform 1 0 1213 0 1 10754
box -255 -1336 255 1336
use sky130_fd_pr__res_xhigh_po_0p35_5BGKTX  XR3 paramcells
timestamp 1718126023
transform 1 0 1213 0 1 8494
box -255 -916 255 916
<< labels >>
flabel metal2 14156 8260 14356 8460 0 FreeSans 256 0 0 0 AOUT
port 6 nsew
flabel metal2 -340 12140 460 12940 0 FreeSans 256 0 0 0 EG_AVDD
port 3 nsew
flabel metal2 -340 1310 460 2110 0 FreeSans 256 0 0 0 EG_AVSS
port 8 nsew
flabel metal2 -340 7370 -140 7570 0 FreeSans 256 0 0 0 XIN
port 4 nsew
flabel metal2 -340 5130 -140 5330 0 FreeSans 256 0 0 0 XOUT
port 1 nsew
flabel metal2 13560 12140 14360 12940 0 FreeSans 256 0 0 0 SG_AVDD
port 2 nsew
flabel metal2 13566 -2990 14366 -2190 0 FreeSans 256 0 0 0 SG_AVSS
port 7 nsew
flabel metal1 9570 -3230 9770 -3030 0 FreeSans 256 0 0 0 EG_IBIAS
port 5 nsew
<< end >>
