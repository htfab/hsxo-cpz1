magic
tech sky130A
magscale 1 2
timestamp 1712819469
<< pwell >>
rect -2727 -3458 2727 3458
<< mvnmos >>
rect -2499 -3200 -2399 3200
rect -2341 -3200 -2241 3200
rect -2183 -3200 -2083 3200
rect -2025 -3200 -1925 3200
rect -1867 -3200 -1767 3200
rect -1709 -3200 -1609 3200
rect -1551 -3200 -1451 3200
rect -1393 -3200 -1293 3200
rect -1235 -3200 -1135 3200
rect -1077 -3200 -977 3200
rect -919 -3200 -819 3200
rect -761 -3200 -661 3200
rect -603 -3200 -503 3200
rect -445 -3200 -345 3200
rect -287 -3200 -187 3200
rect -129 -3200 -29 3200
rect 29 -3200 129 3200
rect 187 -3200 287 3200
rect 345 -3200 445 3200
rect 503 -3200 603 3200
rect 661 -3200 761 3200
rect 819 -3200 919 3200
rect 977 -3200 1077 3200
rect 1135 -3200 1235 3200
rect 1293 -3200 1393 3200
rect 1451 -3200 1551 3200
rect 1609 -3200 1709 3200
rect 1767 -3200 1867 3200
rect 1925 -3200 2025 3200
rect 2083 -3200 2183 3200
rect 2241 -3200 2341 3200
rect 2399 -3200 2499 3200
<< mvndiff >>
rect -2557 3188 -2499 3200
rect -2557 -3188 -2545 3188
rect -2511 -3188 -2499 3188
rect -2557 -3200 -2499 -3188
rect -2399 3188 -2341 3200
rect -2399 -3188 -2387 3188
rect -2353 -3188 -2341 3188
rect -2399 -3200 -2341 -3188
rect -2241 3188 -2183 3200
rect -2241 -3188 -2229 3188
rect -2195 -3188 -2183 3188
rect -2241 -3200 -2183 -3188
rect -2083 3188 -2025 3200
rect -2083 -3188 -2071 3188
rect -2037 -3188 -2025 3188
rect -2083 -3200 -2025 -3188
rect -1925 3188 -1867 3200
rect -1925 -3188 -1913 3188
rect -1879 -3188 -1867 3188
rect -1925 -3200 -1867 -3188
rect -1767 3188 -1709 3200
rect -1767 -3188 -1755 3188
rect -1721 -3188 -1709 3188
rect -1767 -3200 -1709 -3188
rect -1609 3188 -1551 3200
rect -1609 -3188 -1597 3188
rect -1563 -3188 -1551 3188
rect -1609 -3200 -1551 -3188
rect -1451 3188 -1393 3200
rect -1451 -3188 -1439 3188
rect -1405 -3188 -1393 3188
rect -1451 -3200 -1393 -3188
rect -1293 3188 -1235 3200
rect -1293 -3188 -1281 3188
rect -1247 -3188 -1235 3188
rect -1293 -3200 -1235 -3188
rect -1135 3188 -1077 3200
rect -1135 -3188 -1123 3188
rect -1089 -3188 -1077 3188
rect -1135 -3200 -1077 -3188
rect -977 3188 -919 3200
rect -977 -3188 -965 3188
rect -931 -3188 -919 3188
rect -977 -3200 -919 -3188
rect -819 3188 -761 3200
rect -819 -3188 -807 3188
rect -773 -3188 -761 3188
rect -819 -3200 -761 -3188
rect -661 3188 -603 3200
rect -661 -3188 -649 3188
rect -615 -3188 -603 3188
rect -661 -3200 -603 -3188
rect -503 3188 -445 3200
rect -503 -3188 -491 3188
rect -457 -3188 -445 3188
rect -503 -3200 -445 -3188
rect -345 3188 -287 3200
rect -345 -3188 -333 3188
rect -299 -3188 -287 3188
rect -345 -3200 -287 -3188
rect -187 3188 -129 3200
rect -187 -3188 -175 3188
rect -141 -3188 -129 3188
rect -187 -3200 -129 -3188
rect -29 3188 29 3200
rect -29 -3188 -17 3188
rect 17 -3188 29 3188
rect -29 -3200 29 -3188
rect 129 3188 187 3200
rect 129 -3188 141 3188
rect 175 -3188 187 3188
rect 129 -3200 187 -3188
rect 287 3188 345 3200
rect 287 -3188 299 3188
rect 333 -3188 345 3188
rect 287 -3200 345 -3188
rect 445 3188 503 3200
rect 445 -3188 457 3188
rect 491 -3188 503 3188
rect 445 -3200 503 -3188
rect 603 3188 661 3200
rect 603 -3188 615 3188
rect 649 -3188 661 3188
rect 603 -3200 661 -3188
rect 761 3188 819 3200
rect 761 -3188 773 3188
rect 807 -3188 819 3188
rect 761 -3200 819 -3188
rect 919 3188 977 3200
rect 919 -3188 931 3188
rect 965 -3188 977 3188
rect 919 -3200 977 -3188
rect 1077 3188 1135 3200
rect 1077 -3188 1089 3188
rect 1123 -3188 1135 3188
rect 1077 -3200 1135 -3188
rect 1235 3188 1293 3200
rect 1235 -3188 1247 3188
rect 1281 -3188 1293 3188
rect 1235 -3200 1293 -3188
rect 1393 3188 1451 3200
rect 1393 -3188 1405 3188
rect 1439 -3188 1451 3188
rect 1393 -3200 1451 -3188
rect 1551 3188 1609 3200
rect 1551 -3188 1563 3188
rect 1597 -3188 1609 3188
rect 1551 -3200 1609 -3188
rect 1709 3188 1767 3200
rect 1709 -3188 1721 3188
rect 1755 -3188 1767 3188
rect 1709 -3200 1767 -3188
rect 1867 3188 1925 3200
rect 1867 -3188 1879 3188
rect 1913 -3188 1925 3188
rect 1867 -3200 1925 -3188
rect 2025 3188 2083 3200
rect 2025 -3188 2037 3188
rect 2071 -3188 2083 3188
rect 2025 -3200 2083 -3188
rect 2183 3188 2241 3200
rect 2183 -3188 2195 3188
rect 2229 -3188 2241 3188
rect 2183 -3200 2241 -3188
rect 2341 3188 2399 3200
rect 2341 -3188 2353 3188
rect 2387 -3188 2399 3188
rect 2341 -3200 2399 -3188
rect 2499 3188 2557 3200
rect 2499 -3188 2511 3188
rect 2545 -3188 2557 3188
rect 2499 -3200 2557 -3188
<< mvndiffc >>
rect -2545 -3188 -2511 3188
rect -2387 -3188 -2353 3188
rect -2229 -3188 -2195 3188
rect -2071 -3188 -2037 3188
rect -1913 -3188 -1879 3188
rect -1755 -3188 -1721 3188
rect -1597 -3188 -1563 3188
rect -1439 -3188 -1405 3188
rect -1281 -3188 -1247 3188
rect -1123 -3188 -1089 3188
rect -965 -3188 -931 3188
rect -807 -3188 -773 3188
rect -649 -3188 -615 3188
rect -491 -3188 -457 3188
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
rect 457 -3188 491 3188
rect 615 -3188 649 3188
rect 773 -3188 807 3188
rect 931 -3188 965 3188
rect 1089 -3188 1123 3188
rect 1247 -3188 1281 3188
rect 1405 -3188 1439 3188
rect 1563 -3188 1597 3188
rect 1721 -3188 1755 3188
rect 1879 -3188 1913 3188
rect 2037 -3188 2071 3188
rect 2195 -3188 2229 3188
rect 2353 -3188 2387 3188
rect 2511 -3188 2545 3188
<< mvpsubdiff >>
rect -2691 3410 2691 3422
rect -2691 3376 -2583 3410
rect 2583 3376 2691 3410
rect -2691 3364 2691 3376
rect -2691 3314 -2633 3364
rect -2691 -3314 -2679 3314
rect -2645 -3314 -2633 3314
rect 2633 3314 2691 3364
rect -2691 -3364 -2633 -3314
rect 2633 -3314 2645 3314
rect 2679 -3314 2691 3314
rect 2633 -3364 2691 -3314
rect -2691 -3376 2691 -3364
rect -2691 -3410 -2583 -3376
rect 2583 -3410 2691 -3376
rect -2691 -3422 2691 -3410
<< mvpsubdiffcont >>
rect -2583 3376 2583 3410
rect -2679 -3314 -2645 3314
rect 2645 -3314 2679 3314
rect -2583 -3410 2583 -3376
<< poly >>
rect -2499 3272 -2399 3288
rect -2499 3238 -2483 3272
rect -2415 3238 -2399 3272
rect -2499 3200 -2399 3238
rect -2341 3272 -2241 3288
rect -2341 3238 -2325 3272
rect -2257 3238 -2241 3272
rect -2341 3200 -2241 3238
rect -2183 3272 -2083 3288
rect -2183 3238 -2167 3272
rect -2099 3238 -2083 3272
rect -2183 3200 -2083 3238
rect -2025 3272 -1925 3288
rect -2025 3238 -2009 3272
rect -1941 3238 -1925 3272
rect -2025 3200 -1925 3238
rect -1867 3272 -1767 3288
rect -1867 3238 -1851 3272
rect -1783 3238 -1767 3272
rect -1867 3200 -1767 3238
rect -1709 3272 -1609 3288
rect -1709 3238 -1693 3272
rect -1625 3238 -1609 3272
rect -1709 3200 -1609 3238
rect -1551 3272 -1451 3288
rect -1551 3238 -1535 3272
rect -1467 3238 -1451 3272
rect -1551 3200 -1451 3238
rect -1393 3272 -1293 3288
rect -1393 3238 -1377 3272
rect -1309 3238 -1293 3272
rect -1393 3200 -1293 3238
rect -1235 3272 -1135 3288
rect -1235 3238 -1219 3272
rect -1151 3238 -1135 3272
rect -1235 3200 -1135 3238
rect -1077 3272 -977 3288
rect -1077 3238 -1061 3272
rect -993 3238 -977 3272
rect -1077 3200 -977 3238
rect -919 3272 -819 3288
rect -919 3238 -903 3272
rect -835 3238 -819 3272
rect -919 3200 -819 3238
rect -761 3272 -661 3288
rect -761 3238 -745 3272
rect -677 3238 -661 3272
rect -761 3200 -661 3238
rect -603 3272 -503 3288
rect -603 3238 -587 3272
rect -519 3238 -503 3272
rect -603 3200 -503 3238
rect -445 3272 -345 3288
rect -445 3238 -429 3272
rect -361 3238 -345 3272
rect -445 3200 -345 3238
rect -287 3272 -187 3288
rect -287 3238 -271 3272
rect -203 3238 -187 3272
rect -287 3200 -187 3238
rect -129 3272 -29 3288
rect -129 3238 -113 3272
rect -45 3238 -29 3272
rect -129 3200 -29 3238
rect 29 3272 129 3288
rect 29 3238 45 3272
rect 113 3238 129 3272
rect 29 3200 129 3238
rect 187 3272 287 3288
rect 187 3238 203 3272
rect 271 3238 287 3272
rect 187 3200 287 3238
rect 345 3272 445 3288
rect 345 3238 361 3272
rect 429 3238 445 3272
rect 345 3200 445 3238
rect 503 3272 603 3288
rect 503 3238 519 3272
rect 587 3238 603 3272
rect 503 3200 603 3238
rect 661 3272 761 3288
rect 661 3238 677 3272
rect 745 3238 761 3272
rect 661 3200 761 3238
rect 819 3272 919 3288
rect 819 3238 835 3272
rect 903 3238 919 3272
rect 819 3200 919 3238
rect 977 3272 1077 3288
rect 977 3238 993 3272
rect 1061 3238 1077 3272
rect 977 3200 1077 3238
rect 1135 3272 1235 3288
rect 1135 3238 1151 3272
rect 1219 3238 1235 3272
rect 1135 3200 1235 3238
rect 1293 3272 1393 3288
rect 1293 3238 1309 3272
rect 1377 3238 1393 3272
rect 1293 3200 1393 3238
rect 1451 3272 1551 3288
rect 1451 3238 1467 3272
rect 1535 3238 1551 3272
rect 1451 3200 1551 3238
rect 1609 3272 1709 3288
rect 1609 3238 1625 3272
rect 1693 3238 1709 3272
rect 1609 3200 1709 3238
rect 1767 3272 1867 3288
rect 1767 3238 1783 3272
rect 1851 3238 1867 3272
rect 1767 3200 1867 3238
rect 1925 3272 2025 3288
rect 1925 3238 1941 3272
rect 2009 3238 2025 3272
rect 1925 3200 2025 3238
rect 2083 3272 2183 3288
rect 2083 3238 2099 3272
rect 2167 3238 2183 3272
rect 2083 3200 2183 3238
rect 2241 3272 2341 3288
rect 2241 3238 2257 3272
rect 2325 3238 2341 3272
rect 2241 3200 2341 3238
rect 2399 3272 2499 3288
rect 2399 3238 2415 3272
rect 2483 3238 2499 3272
rect 2399 3200 2499 3238
rect -2499 -3238 -2399 -3200
rect -2499 -3272 -2483 -3238
rect -2415 -3272 -2399 -3238
rect -2499 -3288 -2399 -3272
rect -2341 -3238 -2241 -3200
rect -2341 -3272 -2325 -3238
rect -2257 -3272 -2241 -3238
rect -2341 -3288 -2241 -3272
rect -2183 -3238 -2083 -3200
rect -2183 -3272 -2167 -3238
rect -2099 -3272 -2083 -3238
rect -2183 -3288 -2083 -3272
rect -2025 -3238 -1925 -3200
rect -2025 -3272 -2009 -3238
rect -1941 -3272 -1925 -3238
rect -2025 -3288 -1925 -3272
rect -1867 -3238 -1767 -3200
rect -1867 -3272 -1851 -3238
rect -1783 -3272 -1767 -3238
rect -1867 -3288 -1767 -3272
rect -1709 -3238 -1609 -3200
rect -1709 -3272 -1693 -3238
rect -1625 -3272 -1609 -3238
rect -1709 -3288 -1609 -3272
rect -1551 -3238 -1451 -3200
rect -1551 -3272 -1535 -3238
rect -1467 -3272 -1451 -3238
rect -1551 -3288 -1451 -3272
rect -1393 -3238 -1293 -3200
rect -1393 -3272 -1377 -3238
rect -1309 -3272 -1293 -3238
rect -1393 -3288 -1293 -3272
rect -1235 -3238 -1135 -3200
rect -1235 -3272 -1219 -3238
rect -1151 -3272 -1135 -3238
rect -1235 -3288 -1135 -3272
rect -1077 -3238 -977 -3200
rect -1077 -3272 -1061 -3238
rect -993 -3272 -977 -3238
rect -1077 -3288 -977 -3272
rect -919 -3238 -819 -3200
rect -919 -3272 -903 -3238
rect -835 -3272 -819 -3238
rect -919 -3288 -819 -3272
rect -761 -3238 -661 -3200
rect -761 -3272 -745 -3238
rect -677 -3272 -661 -3238
rect -761 -3288 -661 -3272
rect -603 -3238 -503 -3200
rect -603 -3272 -587 -3238
rect -519 -3272 -503 -3238
rect -603 -3288 -503 -3272
rect -445 -3238 -345 -3200
rect -445 -3272 -429 -3238
rect -361 -3272 -345 -3238
rect -445 -3288 -345 -3272
rect -287 -3238 -187 -3200
rect -287 -3272 -271 -3238
rect -203 -3272 -187 -3238
rect -287 -3288 -187 -3272
rect -129 -3238 -29 -3200
rect -129 -3272 -113 -3238
rect -45 -3272 -29 -3238
rect -129 -3288 -29 -3272
rect 29 -3238 129 -3200
rect 29 -3272 45 -3238
rect 113 -3272 129 -3238
rect 29 -3288 129 -3272
rect 187 -3238 287 -3200
rect 187 -3272 203 -3238
rect 271 -3272 287 -3238
rect 187 -3288 287 -3272
rect 345 -3238 445 -3200
rect 345 -3272 361 -3238
rect 429 -3272 445 -3238
rect 345 -3288 445 -3272
rect 503 -3238 603 -3200
rect 503 -3272 519 -3238
rect 587 -3272 603 -3238
rect 503 -3288 603 -3272
rect 661 -3238 761 -3200
rect 661 -3272 677 -3238
rect 745 -3272 761 -3238
rect 661 -3288 761 -3272
rect 819 -3238 919 -3200
rect 819 -3272 835 -3238
rect 903 -3272 919 -3238
rect 819 -3288 919 -3272
rect 977 -3238 1077 -3200
rect 977 -3272 993 -3238
rect 1061 -3272 1077 -3238
rect 977 -3288 1077 -3272
rect 1135 -3238 1235 -3200
rect 1135 -3272 1151 -3238
rect 1219 -3272 1235 -3238
rect 1135 -3288 1235 -3272
rect 1293 -3238 1393 -3200
rect 1293 -3272 1309 -3238
rect 1377 -3272 1393 -3238
rect 1293 -3288 1393 -3272
rect 1451 -3238 1551 -3200
rect 1451 -3272 1467 -3238
rect 1535 -3272 1551 -3238
rect 1451 -3288 1551 -3272
rect 1609 -3238 1709 -3200
rect 1609 -3272 1625 -3238
rect 1693 -3272 1709 -3238
rect 1609 -3288 1709 -3272
rect 1767 -3238 1867 -3200
rect 1767 -3272 1783 -3238
rect 1851 -3272 1867 -3238
rect 1767 -3288 1867 -3272
rect 1925 -3238 2025 -3200
rect 1925 -3272 1941 -3238
rect 2009 -3272 2025 -3238
rect 1925 -3288 2025 -3272
rect 2083 -3238 2183 -3200
rect 2083 -3272 2099 -3238
rect 2167 -3272 2183 -3238
rect 2083 -3288 2183 -3272
rect 2241 -3238 2341 -3200
rect 2241 -3272 2257 -3238
rect 2325 -3272 2341 -3238
rect 2241 -3288 2341 -3272
rect 2399 -3238 2499 -3200
rect 2399 -3272 2415 -3238
rect 2483 -3272 2499 -3238
rect 2399 -3288 2499 -3272
<< polycont >>
rect -2483 3238 -2415 3272
rect -2325 3238 -2257 3272
rect -2167 3238 -2099 3272
rect -2009 3238 -1941 3272
rect -1851 3238 -1783 3272
rect -1693 3238 -1625 3272
rect -1535 3238 -1467 3272
rect -1377 3238 -1309 3272
rect -1219 3238 -1151 3272
rect -1061 3238 -993 3272
rect -903 3238 -835 3272
rect -745 3238 -677 3272
rect -587 3238 -519 3272
rect -429 3238 -361 3272
rect -271 3238 -203 3272
rect -113 3238 -45 3272
rect 45 3238 113 3272
rect 203 3238 271 3272
rect 361 3238 429 3272
rect 519 3238 587 3272
rect 677 3238 745 3272
rect 835 3238 903 3272
rect 993 3238 1061 3272
rect 1151 3238 1219 3272
rect 1309 3238 1377 3272
rect 1467 3238 1535 3272
rect 1625 3238 1693 3272
rect 1783 3238 1851 3272
rect 1941 3238 2009 3272
rect 2099 3238 2167 3272
rect 2257 3238 2325 3272
rect 2415 3238 2483 3272
rect -2483 -3272 -2415 -3238
rect -2325 -3272 -2257 -3238
rect -2167 -3272 -2099 -3238
rect -2009 -3272 -1941 -3238
rect -1851 -3272 -1783 -3238
rect -1693 -3272 -1625 -3238
rect -1535 -3272 -1467 -3238
rect -1377 -3272 -1309 -3238
rect -1219 -3272 -1151 -3238
rect -1061 -3272 -993 -3238
rect -903 -3272 -835 -3238
rect -745 -3272 -677 -3238
rect -587 -3272 -519 -3238
rect -429 -3272 -361 -3238
rect -271 -3272 -203 -3238
rect -113 -3272 -45 -3238
rect 45 -3272 113 -3238
rect 203 -3272 271 -3238
rect 361 -3272 429 -3238
rect 519 -3272 587 -3238
rect 677 -3272 745 -3238
rect 835 -3272 903 -3238
rect 993 -3272 1061 -3238
rect 1151 -3272 1219 -3238
rect 1309 -3272 1377 -3238
rect 1467 -3272 1535 -3238
rect 1625 -3272 1693 -3238
rect 1783 -3272 1851 -3238
rect 1941 -3272 2009 -3238
rect 2099 -3272 2167 -3238
rect 2257 -3272 2325 -3238
rect 2415 -3272 2483 -3238
<< locali >>
rect -2679 3376 -2583 3410
rect 2583 3376 2679 3410
rect -2679 3314 -2645 3376
rect 2645 3314 2679 3376
rect -2499 3238 -2483 3272
rect -2415 3238 -2399 3272
rect -2341 3238 -2325 3272
rect -2257 3238 -2241 3272
rect -2183 3238 -2167 3272
rect -2099 3238 -2083 3272
rect -2025 3238 -2009 3272
rect -1941 3238 -1925 3272
rect -1867 3238 -1851 3272
rect -1783 3238 -1767 3272
rect -1709 3238 -1693 3272
rect -1625 3238 -1609 3272
rect -1551 3238 -1535 3272
rect -1467 3238 -1451 3272
rect -1393 3238 -1377 3272
rect -1309 3238 -1293 3272
rect -1235 3238 -1219 3272
rect -1151 3238 -1135 3272
rect -1077 3238 -1061 3272
rect -993 3238 -977 3272
rect -919 3238 -903 3272
rect -835 3238 -819 3272
rect -761 3238 -745 3272
rect -677 3238 -661 3272
rect -603 3238 -587 3272
rect -519 3238 -503 3272
rect -445 3238 -429 3272
rect -361 3238 -345 3272
rect -287 3238 -271 3272
rect -203 3238 -187 3272
rect -129 3238 -113 3272
rect -45 3238 -29 3272
rect 29 3238 45 3272
rect 113 3238 129 3272
rect 187 3238 203 3272
rect 271 3238 287 3272
rect 345 3238 361 3272
rect 429 3238 445 3272
rect 503 3238 519 3272
rect 587 3238 603 3272
rect 661 3238 677 3272
rect 745 3238 761 3272
rect 819 3238 835 3272
rect 903 3238 919 3272
rect 977 3238 993 3272
rect 1061 3238 1077 3272
rect 1135 3238 1151 3272
rect 1219 3238 1235 3272
rect 1293 3238 1309 3272
rect 1377 3238 1393 3272
rect 1451 3238 1467 3272
rect 1535 3238 1551 3272
rect 1609 3238 1625 3272
rect 1693 3238 1709 3272
rect 1767 3238 1783 3272
rect 1851 3238 1867 3272
rect 1925 3238 1941 3272
rect 2009 3238 2025 3272
rect 2083 3238 2099 3272
rect 2167 3238 2183 3272
rect 2241 3238 2257 3272
rect 2325 3238 2341 3272
rect 2399 3238 2415 3272
rect 2483 3238 2499 3272
rect -2545 3188 -2511 3204
rect -2545 -3204 -2511 -3188
rect -2387 3188 -2353 3204
rect -2387 -3204 -2353 -3188
rect -2229 3188 -2195 3204
rect -2229 -3204 -2195 -3188
rect -2071 3188 -2037 3204
rect -2071 -3204 -2037 -3188
rect -1913 3188 -1879 3204
rect -1913 -3204 -1879 -3188
rect -1755 3188 -1721 3204
rect -1755 -3204 -1721 -3188
rect -1597 3188 -1563 3204
rect -1597 -3204 -1563 -3188
rect -1439 3188 -1405 3204
rect -1439 -3204 -1405 -3188
rect -1281 3188 -1247 3204
rect -1281 -3204 -1247 -3188
rect -1123 3188 -1089 3204
rect -1123 -3204 -1089 -3188
rect -965 3188 -931 3204
rect -965 -3204 -931 -3188
rect -807 3188 -773 3204
rect -807 -3204 -773 -3188
rect -649 3188 -615 3204
rect -649 -3204 -615 -3188
rect -491 3188 -457 3204
rect -491 -3204 -457 -3188
rect -333 3188 -299 3204
rect -333 -3204 -299 -3188
rect -175 3188 -141 3204
rect -175 -3204 -141 -3188
rect -17 3188 17 3204
rect -17 -3204 17 -3188
rect 141 3188 175 3204
rect 141 -3204 175 -3188
rect 299 3188 333 3204
rect 299 -3204 333 -3188
rect 457 3188 491 3204
rect 457 -3204 491 -3188
rect 615 3188 649 3204
rect 615 -3204 649 -3188
rect 773 3188 807 3204
rect 773 -3204 807 -3188
rect 931 3188 965 3204
rect 931 -3204 965 -3188
rect 1089 3188 1123 3204
rect 1089 -3204 1123 -3188
rect 1247 3188 1281 3204
rect 1247 -3204 1281 -3188
rect 1405 3188 1439 3204
rect 1405 -3204 1439 -3188
rect 1563 3188 1597 3204
rect 1563 -3204 1597 -3188
rect 1721 3188 1755 3204
rect 1721 -3204 1755 -3188
rect 1879 3188 1913 3204
rect 1879 -3204 1913 -3188
rect 2037 3188 2071 3204
rect 2037 -3204 2071 -3188
rect 2195 3188 2229 3204
rect 2195 -3204 2229 -3188
rect 2353 3188 2387 3204
rect 2353 -3204 2387 -3188
rect 2511 3188 2545 3204
rect 2511 -3204 2545 -3188
rect -2499 -3272 -2483 -3238
rect -2415 -3272 -2399 -3238
rect -2341 -3272 -2325 -3238
rect -2257 -3272 -2241 -3238
rect -2183 -3272 -2167 -3238
rect -2099 -3272 -2083 -3238
rect -2025 -3272 -2009 -3238
rect -1941 -3272 -1925 -3238
rect -1867 -3272 -1851 -3238
rect -1783 -3272 -1767 -3238
rect -1709 -3272 -1693 -3238
rect -1625 -3272 -1609 -3238
rect -1551 -3272 -1535 -3238
rect -1467 -3272 -1451 -3238
rect -1393 -3272 -1377 -3238
rect -1309 -3272 -1293 -3238
rect -1235 -3272 -1219 -3238
rect -1151 -3272 -1135 -3238
rect -1077 -3272 -1061 -3238
rect -993 -3272 -977 -3238
rect -919 -3272 -903 -3238
rect -835 -3272 -819 -3238
rect -761 -3272 -745 -3238
rect -677 -3272 -661 -3238
rect -603 -3272 -587 -3238
rect -519 -3272 -503 -3238
rect -445 -3272 -429 -3238
rect -361 -3272 -345 -3238
rect -287 -3272 -271 -3238
rect -203 -3272 -187 -3238
rect -129 -3272 -113 -3238
rect -45 -3272 -29 -3238
rect 29 -3272 45 -3238
rect 113 -3272 129 -3238
rect 187 -3272 203 -3238
rect 271 -3272 287 -3238
rect 345 -3272 361 -3238
rect 429 -3272 445 -3238
rect 503 -3272 519 -3238
rect 587 -3272 603 -3238
rect 661 -3272 677 -3238
rect 745 -3272 761 -3238
rect 819 -3272 835 -3238
rect 903 -3272 919 -3238
rect 977 -3272 993 -3238
rect 1061 -3272 1077 -3238
rect 1135 -3272 1151 -3238
rect 1219 -3272 1235 -3238
rect 1293 -3272 1309 -3238
rect 1377 -3272 1393 -3238
rect 1451 -3272 1467 -3238
rect 1535 -3272 1551 -3238
rect 1609 -3272 1625 -3238
rect 1693 -3272 1709 -3238
rect 1767 -3272 1783 -3238
rect 1851 -3272 1867 -3238
rect 1925 -3272 1941 -3238
rect 2009 -3272 2025 -3238
rect 2083 -3272 2099 -3238
rect 2167 -3272 2183 -3238
rect 2241 -3272 2257 -3238
rect 2325 -3272 2341 -3238
rect 2399 -3272 2415 -3238
rect 2483 -3272 2499 -3238
rect -2679 -3376 -2645 -3314
rect 2645 -3376 2679 -3314
rect -2679 -3410 -2583 -3376
rect 2583 -3410 2679 -3376
<< viali >>
rect -2483 3238 -2415 3272
rect -2325 3238 -2257 3272
rect -2167 3238 -2099 3272
rect -2009 3238 -1941 3272
rect -1851 3238 -1783 3272
rect -1693 3238 -1625 3272
rect -1535 3238 -1467 3272
rect -1377 3238 -1309 3272
rect -1219 3238 -1151 3272
rect -1061 3238 -993 3272
rect -903 3238 -835 3272
rect -745 3238 -677 3272
rect -587 3238 -519 3272
rect -429 3238 -361 3272
rect -271 3238 -203 3272
rect -113 3238 -45 3272
rect 45 3238 113 3272
rect 203 3238 271 3272
rect 361 3238 429 3272
rect 519 3238 587 3272
rect 677 3238 745 3272
rect 835 3238 903 3272
rect 993 3238 1061 3272
rect 1151 3238 1219 3272
rect 1309 3238 1377 3272
rect 1467 3238 1535 3272
rect 1625 3238 1693 3272
rect 1783 3238 1851 3272
rect 1941 3238 2009 3272
rect 2099 3238 2167 3272
rect 2257 3238 2325 3272
rect 2415 3238 2483 3272
rect -2545 -3188 -2511 3188
rect -2387 -3188 -2353 3188
rect -2229 -3188 -2195 3188
rect -2071 -3188 -2037 3188
rect -1913 -3188 -1879 3188
rect -1755 -3188 -1721 3188
rect -1597 -3188 -1563 3188
rect -1439 -3188 -1405 3188
rect -1281 -3188 -1247 3188
rect -1123 -3188 -1089 3188
rect -965 -3188 -931 3188
rect -807 -3188 -773 3188
rect -649 -3188 -615 3188
rect -491 -3188 -457 3188
rect -333 -3188 -299 3188
rect -175 -3188 -141 3188
rect -17 -3188 17 3188
rect 141 -3188 175 3188
rect 299 -3188 333 3188
rect 457 -3188 491 3188
rect 615 -3188 649 3188
rect 773 -3188 807 3188
rect 931 -3188 965 3188
rect 1089 -3188 1123 3188
rect 1247 -3188 1281 3188
rect 1405 -3188 1439 3188
rect 1563 -3188 1597 3188
rect 1721 -3188 1755 3188
rect 1879 -3188 1913 3188
rect 2037 -3188 2071 3188
rect 2195 -3188 2229 3188
rect 2353 -3188 2387 3188
rect 2511 -3188 2545 3188
rect -2483 -3272 -2415 -3238
rect -2325 -3272 -2257 -3238
rect -2167 -3272 -2099 -3238
rect -2009 -3272 -1941 -3238
rect -1851 -3272 -1783 -3238
rect -1693 -3272 -1625 -3238
rect -1535 -3272 -1467 -3238
rect -1377 -3272 -1309 -3238
rect -1219 -3272 -1151 -3238
rect -1061 -3272 -993 -3238
rect -903 -3272 -835 -3238
rect -745 -3272 -677 -3238
rect -587 -3272 -519 -3238
rect -429 -3272 -361 -3238
rect -271 -3272 -203 -3238
rect -113 -3272 -45 -3238
rect 45 -3272 113 -3238
rect 203 -3272 271 -3238
rect 361 -3272 429 -3238
rect 519 -3272 587 -3238
rect 677 -3272 745 -3238
rect 835 -3272 903 -3238
rect 993 -3272 1061 -3238
rect 1151 -3272 1219 -3238
rect 1309 -3272 1377 -3238
rect 1467 -3272 1535 -3238
rect 1625 -3272 1693 -3238
rect 1783 -3272 1851 -3238
rect 1941 -3272 2009 -3238
rect 2099 -3272 2167 -3238
rect 2257 -3272 2325 -3238
rect 2415 -3272 2483 -3238
<< metal1 >>
rect -2495 3272 -2403 3278
rect -2495 3238 -2483 3272
rect -2415 3238 -2403 3272
rect -2495 3232 -2403 3238
rect -2337 3272 -2245 3278
rect -2337 3238 -2325 3272
rect -2257 3238 -2245 3272
rect -2337 3232 -2245 3238
rect -2179 3272 -2087 3278
rect -2179 3238 -2167 3272
rect -2099 3238 -2087 3272
rect -2179 3232 -2087 3238
rect -2021 3272 -1929 3278
rect -2021 3238 -2009 3272
rect -1941 3238 -1929 3272
rect -2021 3232 -1929 3238
rect -1863 3272 -1771 3278
rect -1863 3238 -1851 3272
rect -1783 3238 -1771 3272
rect -1863 3232 -1771 3238
rect -1705 3272 -1613 3278
rect -1705 3238 -1693 3272
rect -1625 3238 -1613 3272
rect -1705 3232 -1613 3238
rect -1547 3272 -1455 3278
rect -1547 3238 -1535 3272
rect -1467 3238 -1455 3272
rect -1547 3232 -1455 3238
rect -1389 3272 -1297 3278
rect -1389 3238 -1377 3272
rect -1309 3238 -1297 3272
rect -1389 3232 -1297 3238
rect -1231 3272 -1139 3278
rect -1231 3238 -1219 3272
rect -1151 3238 -1139 3272
rect -1231 3232 -1139 3238
rect -1073 3272 -981 3278
rect -1073 3238 -1061 3272
rect -993 3238 -981 3272
rect -1073 3232 -981 3238
rect -915 3272 -823 3278
rect -915 3238 -903 3272
rect -835 3238 -823 3272
rect -915 3232 -823 3238
rect -757 3272 -665 3278
rect -757 3238 -745 3272
rect -677 3238 -665 3272
rect -757 3232 -665 3238
rect -599 3272 -507 3278
rect -599 3238 -587 3272
rect -519 3238 -507 3272
rect -599 3232 -507 3238
rect -441 3272 -349 3278
rect -441 3238 -429 3272
rect -361 3238 -349 3272
rect -441 3232 -349 3238
rect -283 3272 -191 3278
rect -283 3238 -271 3272
rect -203 3238 -191 3272
rect -283 3232 -191 3238
rect -125 3272 -33 3278
rect -125 3238 -113 3272
rect -45 3238 -33 3272
rect -125 3232 -33 3238
rect 33 3272 125 3278
rect 33 3238 45 3272
rect 113 3238 125 3272
rect 33 3232 125 3238
rect 191 3272 283 3278
rect 191 3238 203 3272
rect 271 3238 283 3272
rect 191 3232 283 3238
rect 349 3272 441 3278
rect 349 3238 361 3272
rect 429 3238 441 3272
rect 349 3232 441 3238
rect 507 3272 599 3278
rect 507 3238 519 3272
rect 587 3238 599 3272
rect 507 3232 599 3238
rect 665 3272 757 3278
rect 665 3238 677 3272
rect 745 3238 757 3272
rect 665 3232 757 3238
rect 823 3272 915 3278
rect 823 3238 835 3272
rect 903 3238 915 3272
rect 823 3232 915 3238
rect 981 3272 1073 3278
rect 981 3238 993 3272
rect 1061 3238 1073 3272
rect 981 3232 1073 3238
rect 1139 3272 1231 3278
rect 1139 3238 1151 3272
rect 1219 3238 1231 3272
rect 1139 3232 1231 3238
rect 1297 3272 1389 3278
rect 1297 3238 1309 3272
rect 1377 3238 1389 3272
rect 1297 3232 1389 3238
rect 1455 3272 1547 3278
rect 1455 3238 1467 3272
rect 1535 3238 1547 3272
rect 1455 3232 1547 3238
rect 1613 3272 1705 3278
rect 1613 3238 1625 3272
rect 1693 3238 1705 3272
rect 1613 3232 1705 3238
rect 1771 3272 1863 3278
rect 1771 3238 1783 3272
rect 1851 3238 1863 3272
rect 1771 3232 1863 3238
rect 1929 3272 2021 3278
rect 1929 3238 1941 3272
rect 2009 3238 2021 3272
rect 1929 3232 2021 3238
rect 2087 3272 2179 3278
rect 2087 3238 2099 3272
rect 2167 3238 2179 3272
rect 2087 3232 2179 3238
rect 2245 3272 2337 3278
rect 2245 3238 2257 3272
rect 2325 3238 2337 3272
rect 2245 3232 2337 3238
rect 2403 3272 2495 3278
rect 2403 3238 2415 3272
rect 2483 3238 2495 3272
rect 2403 3232 2495 3238
rect -2551 3188 -2505 3200
rect -2551 -3188 -2545 3188
rect -2511 -3188 -2505 3188
rect -2551 -3200 -2505 -3188
rect -2393 3188 -2347 3200
rect -2393 -3188 -2387 3188
rect -2353 -3188 -2347 3188
rect -2393 -3200 -2347 -3188
rect -2235 3188 -2189 3200
rect -2235 -3188 -2229 3188
rect -2195 -3188 -2189 3188
rect -2235 -3200 -2189 -3188
rect -2077 3188 -2031 3200
rect -2077 -3188 -2071 3188
rect -2037 -3188 -2031 3188
rect -2077 -3200 -2031 -3188
rect -1919 3188 -1873 3200
rect -1919 -3188 -1913 3188
rect -1879 -3188 -1873 3188
rect -1919 -3200 -1873 -3188
rect -1761 3188 -1715 3200
rect -1761 -3188 -1755 3188
rect -1721 -3188 -1715 3188
rect -1761 -3200 -1715 -3188
rect -1603 3188 -1557 3200
rect -1603 -3188 -1597 3188
rect -1563 -3188 -1557 3188
rect -1603 -3200 -1557 -3188
rect -1445 3188 -1399 3200
rect -1445 -3188 -1439 3188
rect -1405 -3188 -1399 3188
rect -1445 -3200 -1399 -3188
rect -1287 3188 -1241 3200
rect -1287 -3188 -1281 3188
rect -1247 -3188 -1241 3188
rect -1287 -3200 -1241 -3188
rect -1129 3188 -1083 3200
rect -1129 -3188 -1123 3188
rect -1089 -3188 -1083 3188
rect -1129 -3200 -1083 -3188
rect -971 3188 -925 3200
rect -971 -3188 -965 3188
rect -931 -3188 -925 3188
rect -971 -3200 -925 -3188
rect -813 3188 -767 3200
rect -813 -3188 -807 3188
rect -773 -3188 -767 3188
rect -813 -3200 -767 -3188
rect -655 3188 -609 3200
rect -655 -3188 -649 3188
rect -615 -3188 -609 3188
rect -655 -3200 -609 -3188
rect -497 3188 -451 3200
rect -497 -3188 -491 3188
rect -457 -3188 -451 3188
rect -497 -3200 -451 -3188
rect -339 3188 -293 3200
rect -339 -3188 -333 3188
rect -299 -3188 -293 3188
rect -339 -3200 -293 -3188
rect -181 3188 -135 3200
rect -181 -3188 -175 3188
rect -141 -3188 -135 3188
rect -181 -3200 -135 -3188
rect -23 3188 23 3200
rect -23 -3188 -17 3188
rect 17 -3188 23 3188
rect -23 -3200 23 -3188
rect 135 3188 181 3200
rect 135 -3188 141 3188
rect 175 -3188 181 3188
rect 135 -3200 181 -3188
rect 293 3188 339 3200
rect 293 -3188 299 3188
rect 333 -3188 339 3188
rect 293 -3200 339 -3188
rect 451 3188 497 3200
rect 451 -3188 457 3188
rect 491 -3188 497 3188
rect 451 -3200 497 -3188
rect 609 3188 655 3200
rect 609 -3188 615 3188
rect 649 -3188 655 3188
rect 609 -3200 655 -3188
rect 767 3188 813 3200
rect 767 -3188 773 3188
rect 807 -3188 813 3188
rect 767 -3200 813 -3188
rect 925 3188 971 3200
rect 925 -3188 931 3188
rect 965 -3188 971 3188
rect 925 -3200 971 -3188
rect 1083 3188 1129 3200
rect 1083 -3188 1089 3188
rect 1123 -3188 1129 3188
rect 1083 -3200 1129 -3188
rect 1241 3188 1287 3200
rect 1241 -3188 1247 3188
rect 1281 -3188 1287 3188
rect 1241 -3200 1287 -3188
rect 1399 3188 1445 3200
rect 1399 -3188 1405 3188
rect 1439 -3188 1445 3188
rect 1399 -3200 1445 -3188
rect 1557 3188 1603 3200
rect 1557 -3188 1563 3188
rect 1597 -3188 1603 3188
rect 1557 -3200 1603 -3188
rect 1715 3188 1761 3200
rect 1715 -3188 1721 3188
rect 1755 -3188 1761 3188
rect 1715 -3200 1761 -3188
rect 1873 3188 1919 3200
rect 1873 -3188 1879 3188
rect 1913 -3188 1919 3188
rect 1873 -3200 1919 -3188
rect 2031 3188 2077 3200
rect 2031 -3188 2037 3188
rect 2071 -3188 2077 3188
rect 2031 -3200 2077 -3188
rect 2189 3188 2235 3200
rect 2189 -3188 2195 3188
rect 2229 -3188 2235 3188
rect 2189 -3200 2235 -3188
rect 2347 3188 2393 3200
rect 2347 -3188 2353 3188
rect 2387 -3188 2393 3188
rect 2347 -3200 2393 -3188
rect 2505 3188 2551 3200
rect 2505 -3188 2511 3188
rect 2545 -3188 2551 3188
rect 2505 -3200 2551 -3188
rect -2495 -3238 -2403 -3232
rect -2495 -3272 -2483 -3238
rect -2415 -3272 -2403 -3238
rect -2495 -3278 -2403 -3272
rect -2337 -3238 -2245 -3232
rect -2337 -3272 -2325 -3238
rect -2257 -3272 -2245 -3238
rect -2337 -3278 -2245 -3272
rect -2179 -3238 -2087 -3232
rect -2179 -3272 -2167 -3238
rect -2099 -3272 -2087 -3238
rect -2179 -3278 -2087 -3272
rect -2021 -3238 -1929 -3232
rect -2021 -3272 -2009 -3238
rect -1941 -3272 -1929 -3238
rect -2021 -3278 -1929 -3272
rect -1863 -3238 -1771 -3232
rect -1863 -3272 -1851 -3238
rect -1783 -3272 -1771 -3238
rect -1863 -3278 -1771 -3272
rect -1705 -3238 -1613 -3232
rect -1705 -3272 -1693 -3238
rect -1625 -3272 -1613 -3238
rect -1705 -3278 -1613 -3272
rect -1547 -3238 -1455 -3232
rect -1547 -3272 -1535 -3238
rect -1467 -3272 -1455 -3238
rect -1547 -3278 -1455 -3272
rect -1389 -3238 -1297 -3232
rect -1389 -3272 -1377 -3238
rect -1309 -3272 -1297 -3238
rect -1389 -3278 -1297 -3272
rect -1231 -3238 -1139 -3232
rect -1231 -3272 -1219 -3238
rect -1151 -3272 -1139 -3238
rect -1231 -3278 -1139 -3272
rect -1073 -3238 -981 -3232
rect -1073 -3272 -1061 -3238
rect -993 -3272 -981 -3238
rect -1073 -3278 -981 -3272
rect -915 -3238 -823 -3232
rect -915 -3272 -903 -3238
rect -835 -3272 -823 -3238
rect -915 -3278 -823 -3272
rect -757 -3238 -665 -3232
rect -757 -3272 -745 -3238
rect -677 -3272 -665 -3238
rect -757 -3278 -665 -3272
rect -599 -3238 -507 -3232
rect -599 -3272 -587 -3238
rect -519 -3272 -507 -3238
rect -599 -3278 -507 -3272
rect -441 -3238 -349 -3232
rect -441 -3272 -429 -3238
rect -361 -3272 -349 -3238
rect -441 -3278 -349 -3272
rect -283 -3238 -191 -3232
rect -283 -3272 -271 -3238
rect -203 -3272 -191 -3238
rect -283 -3278 -191 -3272
rect -125 -3238 -33 -3232
rect -125 -3272 -113 -3238
rect -45 -3272 -33 -3238
rect -125 -3278 -33 -3272
rect 33 -3238 125 -3232
rect 33 -3272 45 -3238
rect 113 -3272 125 -3238
rect 33 -3278 125 -3272
rect 191 -3238 283 -3232
rect 191 -3272 203 -3238
rect 271 -3272 283 -3238
rect 191 -3278 283 -3272
rect 349 -3238 441 -3232
rect 349 -3272 361 -3238
rect 429 -3272 441 -3238
rect 349 -3278 441 -3272
rect 507 -3238 599 -3232
rect 507 -3272 519 -3238
rect 587 -3272 599 -3238
rect 507 -3278 599 -3272
rect 665 -3238 757 -3232
rect 665 -3272 677 -3238
rect 745 -3272 757 -3238
rect 665 -3278 757 -3272
rect 823 -3238 915 -3232
rect 823 -3272 835 -3238
rect 903 -3272 915 -3238
rect 823 -3278 915 -3272
rect 981 -3238 1073 -3232
rect 981 -3272 993 -3238
rect 1061 -3272 1073 -3238
rect 981 -3278 1073 -3272
rect 1139 -3238 1231 -3232
rect 1139 -3272 1151 -3238
rect 1219 -3272 1231 -3238
rect 1139 -3278 1231 -3272
rect 1297 -3238 1389 -3232
rect 1297 -3272 1309 -3238
rect 1377 -3272 1389 -3238
rect 1297 -3278 1389 -3272
rect 1455 -3238 1547 -3232
rect 1455 -3272 1467 -3238
rect 1535 -3272 1547 -3238
rect 1455 -3278 1547 -3272
rect 1613 -3238 1705 -3232
rect 1613 -3272 1625 -3238
rect 1693 -3272 1705 -3238
rect 1613 -3278 1705 -3272
rect 1771 -3238 1863 -3232
rect 1771 -3272 1783 -3238
rect 1851 -3272 1863 -3238
rect 1771 -3278 1863 -3272
rect 1929 -3238 2021 -3232
rect 1929 -3272 1941 -3238
rect 2009 -3272 2021 -3238
rect 1929 -3278 2021 -3272
rect 2087 -3238 2179 -3232
rect 2087 -3272 2099 -3238
rect 2167 -3272 2179 -3238
rect 2087 -3278 2179 -3272
rect 2245 -3238 2337 -3232
rect 2245 -3272 2257 -3238
rect 2325 -3272 2337 -3238
rect 2245 -3278 2337 -3272
rect 2403 -3238 2495 -3232
rect 2403 -3272 2415 -3238
rect 2483 -3272 2495 -3238
rect 2403 -3278 2495 -3272
<< properties >>
string FIXED_BBOX -2662 -3393 2662 3393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 0.5 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
