magic
tech sky130A
magscale 1 2
timestamp 1713791295
<< error_p >>
rect -77 481 -19 487
rect 115 481 173 487
rect -77 447 -65 481
rect 115 447 127 481
rect -77 441 -19 447
rect 115 441 173 447
rect -173 -447 -115 -441
rect 19 -447 77 -441
rect -173 -481 -161 -447
rect 19 -481 31 -447
rect -173 -487 -115 -481
rect 19 -487 77 -481
<< nwell >>
rect -359 -619 359 619
<< pmos >>
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
<< pdiff >>
rect -221 388 -159 400
rect -221 -388 -209 388
rect -175 -388 -159 388
rect -221 -400 -159 -388
rect -129 388 -63 400
rect -129 -388 -113 388
rect -79 -388 -63 388
rect -129 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 129 400
rect 63 -388 79 388
rect 113 -388 129 388
rect 63 -400 129 -388
rect 159 388 221 400
rect 159 -388 175 388
rect 209 -388 221 388
rect 159 -400 221 -388
<< pdiffc >>
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
<< nsubdiff >>
rect -323 549 -227 583
rect 227 549 323 583
rect -323 487 -289 549
rect 289 487 323 549
rect -323 -549 -289 -487
rect 289 -549 323 -487
rect -323 -583 -227 -549
rect 227 -583 323 -549
<< nsubdiffcont >>
rect -227 549 227 583
rect -323 -487 -289 487
rect 289 -487 323 487
rect -227 -583 227 -549
<< poly >>
rect -81 481 -15 497
rect -81 447 -65 481
rect -31 447 -15 481
rect -81 431 -15 447
rect 111 481 177 497
rect 111 447 127 481
rect 161 447 177 481
rect 111 431 177 447
rect -159 400 -129 426
rect -63 400 -33 431
rect 33 400 63 426
rect 129 400 159 431
rect -159 -431 -129 -400
rect -63 -426 -33 -400
rect 33 -431 63 -400
rect 129 -426 159 -400
rect -177 -447 -111 -431
rect -177 -481 -161 -447
rect -127 -481 -111 -447
rect -177 -497 -111 -481
rect 15 -447 81 -431
rect 15 -481 31 -447
rect 65 -481 81 -447
rect 15 -497 81 -481
<< polycont >>
rect -65 447 -31 481
rect 127 447 161 481
rect -161 -481 -127 -447
rect 31 -481 65 -447
<< locali >>
rect -323 549 -227 583
rect 227 549 323 583
rect -323 487 -289 549
rect 289 487 323 549
rect -81 447 -65 481
rect -31 447 -15 481
rect 111 447 127 481
rect 161 447 177 481
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect -177 -481 -161 -447
rect -127 -481 -111 -447
rect 15 -481 31 -447
rect 65 -481 81 -447
rect -323 -549 -289 -487
rect 289 -549 323 -487
rect -323 -583 -227 -549
rect 227 -583 323 -549
<< viali >>
rect -65 447 -31 481
rect 127 447 161 481
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect -161 -481 -127 -447
rect 31 -481 65 -447
<< metal1 >>
rect -77 481 -19 487
rect -77 447 -65 481
rect -31 447 -19 481
rect -77 441 -19 447
rect 115 481 173 487
rect 115 447 127 481
rect 161 447 173 481
rect 115 441 173 447
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect -173 -447 -115 -441
rect -173 -481 -161 -447
rect -127 -481 -115 -447
rect -173 -487 -115 -481
rect 19 -447 77 -441
rect 19 -481 31 -447
rect 65 -481 77 -447
rect 19 -487 77 -481
<< properties >>
string FIXED_BBOX -306 -566 306 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
