magic
tech sky130A
magscale 1 2
timestamp 1713249912
<< pwell >>
rect -193 -193 193 193
<< mvpsubdiff >>
rect -157 123 -51 157
rect 51 123 157 157
rect -157 51 -123 123
rect 123 51 157 123
rect -157 -123 -123 -51
rect 123 -123 157 -51
rect -157 -157 -51 -123
rect 51 -157 157 -123
<< mvpsubdiffcont >>
rect -51 123 51 157
rect -157 -51 -123 51
rect 123 -51 157 51
rect -51 -157 51 -123
<< mvndiode >>
rect -45 33 45 45
rect -49 -33 -33 33
rect 33 -33 49 33
rect -45 -45 45 -33
<< mvndiodec >>
rect -33 -33 33 33
<< locali >>
rect -157 123 -51 157
rect 51 123 157 157
rect -157 51 -123 123
rect 123 51 157 123
rect -49 -33 -33 33
rect 33 -33 49 33
rect -157 -123 -123 -51
rect 123 -123 157 -51
rect -157 -157 -51 -123
rect 51 -157 157 -123
<< viali >>
rect -33 -33 33 33
<< metal1 >>
rect -45 33 45 39
rect -45 -33 -33 33
rect 33 -33 45 33
rect -45 -39 45 -33
<< properties >>
string FIXED_BBOX -130 -130 130 130
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 0.45 l 0.45 area 202.5m peri 1.8 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
