magic
tech sky130A
magscale 1 2
timestamp 1713806792
<< error_s >>
rect 236 12879 256 13084
rect 242 9030 256 12879
rect 244 7942 256 9030
rect 722 8355 734 8989
rect 750 8383 762 9017
rect 722 8191 738 8355
rect 722 8189 734 8191
rect 750 8163 766 8383
rect 750 8161 762 8163
rect 1102 -3914 1128 -3906
rect 1130 -3914 1156 -3878
<< metal1 >>
rect 0 16110 30870 16310
rect 31070 16110 31076 16310
rect 0 602 200 16110
rect 8834 14970 8840 15170
rect 9040 14970 24190 15170
rect 24390 14970 24396 15170
rect 9704 9950 9710 10150
rect 9910 9950 9916 10150
rect 744 9510 750 9710
rect 950 9510 956 9710
rect 364 7042 370 7250
rect 570 7042 576 7250
rect -6 400 0 602
rect 200 400 206 602
rect 370 -6750 570 7042
rect 750 5572 950 9510
rect 8840 7012 9040 7018
rect 9710 7012 9910 9950
rect 9040 6812 9910 7012
rect 8840 6806 9040 6812
rect 8834 6390 8840 6590
rect 9040 6390 9480 6590
rect 8824 6000 8830 6200
rect 9030 6000 9036 6200
rect 744 5372 750 5572
rect 950 5372 956 5572
rect 1124 -348 1130 -148
rect 1330 -348 1336 -148
rect 1130 -6340 1330 -348
rect 8830 -630 9030 6000
rect 8824 -830 8830 -630
rect 9030 -830 9036 -630
rect 9280 -680 9480 6390
rect 9280 -880 9710 -680
rect 9910 -880 9916 -680
rect 30870 -4510 31070 -4504
rect 30870 -6340 31070 -4710
rect 1130 -6540 31070 -6340
rect 370 -6950 19620 -6750
rect 19820 -6950 19826 -6750
<< via1 >>
rect 30870 16110 31070 16310
rect 8840 14970 9040 15170
rect 24190 14970 24390 15170
rect 9710 9950 9910 10150
rect 750 9510 950 9710
rect 370 7042 570 7250
rect 0 400 200 602
rect 8840 6812 9040 7012
rect 8840 6390 9040 6590
rect 8830 6000 9030 6200
rect 750 5372 950 5572
rect 1130 -348 1330 -148
rect 8830 -830 9030 -630
rect 9710 -880 9910 -680
rect 30870 -4710 31070 -4510
rect 19620 -6950 19820 -6750
<< metal2 >>
rect 30870 16310 31070 16316
rect 0 16305 200 16310
rect -4 16115 5 16305
rect 195 16115 204 16305
rect 0 6860 200 16115
rect 370 16110 9480 16310
rect 370 9280 570 16110
rect 8840 15170 9040 15176
rect 1121 11302 1130 11502
rect 1330 11302 1339 11502
rect 750 9710 950 9716
rect 741 9510 750 9710
rect 950 9510 959 9710
rect 750 9504 950 9510
rect 370 9080 950 9280
rect 370 7250 570 7256
rect 361 7050 370 7250
rect 570 7050 579 7250
rect 366 7047 370 7050
rect 570 7047 574 7050
rect 370 7036 570 7042
rect 0 6651 200 6660
rect 750 5977 950 9080
rect 1121 7442 1130 7642
rect 1330 7442 1339 7642
rect 1121 7042 1130 7242
rect 1330 7042 1339 7242
rect 8840 7172 9040 14970
rect 8834 6812 8840 7012
rect 9040 6812 9046 7012
rect 8840 6590 9040 6596
rect 8840 6384 9040 6390
rect 8830 6200 9030 6206
rect 8830 5994 9030 6000
rect 750 5787 755 5977
rect 945 5787 950 5977
rect 750 5782 950 5787
rect 1121 5782 1130 5982
rect 1330 5782 1339 5982
rect 755 5778 945 5782
rect 750 5572 950 5578
rect 950 5372 1330 5572
rect 9280 5380 9480 16110
rect 25870 16050 26070 16059
rect 30870 15900 31070 16110
rect 24190 15170 24390 15176
rect 9710 10150 9910 10156
rect 24190 9950 24390 14970
rect 9710 9944 9910 9950
rect 25870 6270 26070 15850
rect 24200 6070 26070 6270
rect 750 5366 950 5372
rect 9280 5180 9910 5380
rect 9271 2940 9280 3140
rect 9480 2940 9910 3140
rect 1121 1872 1130 2072
rect 1330 1872 1339 2072
rect 730 1550 930 1559
rect 0 602 200 608
rect -9 400 0 600
rect 200 400 209 600
rect 0 394 200 400
rect 730 237 930 1350
rect 1121 742 1130 942
rect 1330 742 1339 942
rect 1121 402 1130 602
rect 1330 402 1339 602
rect 730 47 735 237
rect 925 47 930 237
rect 730 42 930 47
rect 1121 42 1130 242
rect 1330 42 1339 242
rect 27640 100 27980 300
rect 735 38 925 42
rect 1130 -148 1330 -142
rect 1130 -354 1330 -348
rect 8830 -148 9030 -139
rect 8830 -357 9030 -348
rect 1121 -688 1130 -488
rect 1330 -688 1339 -488
rect 8830 -630 9030 -624
rect 8830 -6340 9030 -830
rect 9710 -680 9910 -674
rect 9710 -886 9910 -880
rect 19155 -6340 19345 -6336
rect 8830 -6345 19350 -6340
rect 8830 -6535 19155 -6345
rect 19345 -6535 19350 -6345
rect 8830 -6540 19350 -6535
rect 19155 -6544 19345 -6540
rect 19620 -6750 19820 -5920
rect 24210 -6340 24410 -4320
rect 27640 -4510 27840 100
rect 30864 -4710 30870 -4510
rect 31070 -4710 31076 -4510
rect 27640 -4719 27840 -4710
rect 20091 -6540 20100 -6340
rect 20300 -6540 24410 -6340
rect 31540 -6750 31740 300
rect 31531 -6950 31540 -6750
rect 31740 -6950 31749 -6750
rect 19620 -6956 19820 -6950
<< via2 >>
rect 5 16115 195 16305
rect 1130 11302 1330 11502
rect 750 9510 950 9710
rect 370 7050 570 7250
rect 375 7047 565 7050
rect 0 6660 200 6860
rect 1130 7442 1330 7642
rect 1130 7042 1330 7242
rect 755 5787 945 5977
rect 1130 5782 1330 5982
rect 25870 15850 26070 16050
rect 9280 2940 9480 3140
rect 1130 1872 1330 2072
rect 730 1350 930 1550
rect 0 400 200 600
rect 1130 742 1330 942
rect 1130 402 1330 602
rect 735 47 925 237
rect 1130 42 1330 242
rect 8830 -348 9030 -148
rect 1130 -688 1330 -488
rect 19155 -6535 19345 -6345
rect 27640 -4710 27840 -4510
rect 20100 -6540 20300 -6340
rect 31540 -6950 31740 -6750
<< metal3 >>
rect 0 16305 9480 16310
rect 0 16115 5 16305
rect 195 16115 9480 16305
rect 0 16110 9480 16115
rect 1125 11502 1335 11507
rect -200 11302 1130 11502
rect 1330 11302 1335 11502
rect -200 11300 0 11302
rect 1125 11297 1335 11302
rect 745 9710 955 9715
rect -200 9510 750 9710
rect 950 9510 955 9710
rect 745 9505 955 9510
rect 1125 7642 1335 7647
rect -200 7442 1130 7642
rect 1330 7442 1335 7642
rect -200 7440 0 7442
rect 1125 7437 1335 7442
rect 365 7250 575 7255
rect 365 7050 370 7250
rect 570 7242 575 7250
rect 1125 7242 1335 7247
rect 570 7050 1130 7242
rect 365 7047 375 7050
rect 565 7047 1130 7050
rect 365 7045 1130 7047
rect 370 7042 1130 7045
rect 1330 7042 1335 7242
rect 1125 7037 1335 7042
rect -5 6860 205 6865
rect -200 6660 0 6860
rect 200 6660 205 6860
rect -5 6655 205 6660
rect 1125 5982 1335 5987
rect -200 5977 1130 5982
rect -200 5787 755 5977
rect 945 5787 1130 5977
rect -200 5782 1130 5787
rect 1330 5782 1335 5982
rect -200 5780 0 5782
rect 1125 5777 1335 5782
rect 9280 3145 9480 16110
rect 25865 16050 26075 16055
rect 25865 16045 25870 16050
rect 26070 16045 26075 16050
rect 25865 15839 26075 15845
rect 9275 3140 9485 3145
rect 9275 2940 9280 3140
rect 9480 2940 9485 3140
rect 9275 2935 9485 2940
rect 1125 2072 1335 2077
rect -200 1872 1130 2072
rect 1330 1872 1335 2072
rect -200 1870 0 1872
rect 1125 1867 1335 1872
rect 725 1550 935 1555
rect -200 1350 730 1550
rect 930 1350 935 1550
rect 725 1345 935 1350
rect 1125 942 1335 947
rect -200 742 1130 942
rect 1330 742 1335 942
rect -200 740 0 742
rect 1125 737 1335 742
rect -5 602 205 605
rect 1125 602 1335 607
rect -5 600 1130 602
rect -5 400 0 600
rect 200 402 1130 600
rect 1330 402 1335 602
rect 200 400 205 402
rect -5 395 205 400
rect 1125 397 1335 402
rect 1125 242 1335 247
rect 730 237 1130 242
rect 730 47 735 237
rect 925 47 1130 237
rect 730 42 1130 47
rect 1330 42 1335 242
rect 1125 37 1335 42
rect 8825 -148 9035 -143
rect 8825 -348 8830 -148
rect 9030 -348 9035 -148
rect 8825 -353 9035 -348
rect 1125 -488 1335 -483
rect -200 -688 1130 -488
rect 1330 -688 1335 -488
rect -200 -690 0 -688
rect 1125 -693 1335 -688
rect 8830 -6750 9030 -353
rect 27635 -4505 27845 -4499
rect 27635 -4710 27640 -4705
rect 27840 -4710 27845 -4705
rect 27635 -4715 27845 -4710
rect 20095 -6340 20305 -6335
rect 19150 -6345 20100 -6340
rect 19150 -6535 19155 -6345
rect 19345 -6535 20100 -6345
rect 19150 -6540 20100 -6535
rect 20300 -6540 20305 -6340
rect 20095 -6545 20305 -6540
rect 31535 -6750 31745 -6745
rect 8830 -6950 31540 -6750
rect 31740 -6950 31950 -6750
rect 31535 -6955 31745 -6950
<< via3 >>
rect 25865 15850 25870 16045
rect 25870 15850 26070 16045
rect 26070 15850 26075 16045
rect 25865 15845 26075 15850
rect 27635 -4510 27845 -4505
rect 27635 -4705 27640 -4510
rect 27640 -4705 27840 -4510
rect 27840 -4705 27845 -4510
<< metal4 >>
rect 25864 16045 26076 16046
rect 25864 15845 25865 16045
rect 26075 15845 26076 16045
rect 25864 15844 26076 15845
rect 25870 -4260 26070 15844
rect 27640 -4504 27840 15660
rect 27634 -4505 27846 -4504
rect 27634 -4705 27635 -4505
rect 27845 -4705 27846 -4505
rect 27634 -4706 27846 -4705
use power_gating  power_gating_0
timestamp 1713806792
transform 1 0 1870 0 1 10256
box -3950 -15179 6766 6365
use schmitt_trigger_pullmid  schmitt_trigger_pullmid_0
timestamp 1713804741
transform 1 0 26390 0 1 -720
box 1390 -3990 5350 16820
use sky130_fd_pr__cap_mim_m3_1_MPZGNS  sky130_fd_pr__cap_mim_m3_1_MPZGNS_0
timestamp 1713804741
transform 1 0 26106 0 1 5700
box -1686 -9960 1686 9960
use vittoz_pierce_osc  vittoz_pierce_osc_0
timestamp 1713804741
transform 1 0 10050 0 1 -2190
box -340 -3940 14370 18841
<< labels >>
flabel metal3 -200 11300 0 11500 0 FreeSans 256 0 0 0 AVDD
port 5 nsew
flabel metal3 -200 9510 0 9710 0 FreeSans 256 0 0 0 AVSS
port 7 nsew
flabel metal3 -200 7440 0 7640 0 FreeSans 256 0 0 0 IBIAS
port 9 nsew
flabel metal3 -200 6660 0 6860 0 FreeSans 256 0 0 0 XOUT
port 0 nsew
flabel metal3 -200 5780 0 5980 0 FreeSans 256 0 0 0 XIN
port 1 nsew
flabel metal3 -200 1870 0 2070 0 FreeSans 256 0 0 0 ENA
port 2 nsew
flabel metal3 -200 1350 0 1550 0 FreeSans 256 0 0 0 STDBY
port 3 nsew
flabel metal3 -200 740 0 940 0 FreeSans 256 0 0 0 DVDD
port 6 nsew
flabel metal3 -200 -690 0 -490 0 FreeSans 256 0 0 0 DVSS
port 8 nsew
flabel metal3 31750 -6950 31950 -6750 0 FreeSans 256 0 0 0 DOUT
port 4 nsew
<< end >>
