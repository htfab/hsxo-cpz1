magic
tech sky130A
magscale 1 2
timestamp 1718126023
<< pwell >>
rect -255 -916 255 916
<< mvpsubdiff >>
rect -189 838 189 850
rect -189 804 -81 838
rect 81 804 189 838
rect -189 792 189 804
rect -189 742 -131 792
rect -189 -742 -177 742
rect -143 -742 -131 742
rect 131 742 189 792
rect -189 -792 -131 -742
rect 131 -742 143 742
rect 177 -742 189 742
rect 131 -792 189 -742
rect -189 -804 189 -792
rect -189 -838 -81 -804
rect 81 -838 189 -804
rect -189 -850 189 -838
<< mvpsubdiffcont >>
rect -81 804 81 838
rect -177 -742 -143 742
rect 143 -742 177 742
rect -81 -838 81 -804
<< xpolycontact >>
rect -35 264 35 696
rect -35 -696 35 -264
<< xpolyres >>
rect -35 -264 35 264
<< locali >>
rect -177 804 -81 838
rect 81 804 177 838
rect -177 742 -143 804
rect 143 742 177 804
rect -177 -804 -143 -742
rect 143 -804 177 -742
rect -177 -838 -81 -804
rect 81 -838 177 -804
<< viali >>
rect -19 281 19 678
rect -19 -678 19 -281
<< metal1 >>
rect -25 678 25 690
rect -25 281 -19 678
rect 19 281 25 678
rect -25 269 25 281
rect -25 -281 25 -269
rect -25 -678 -19 -281
rect 19 -678 25 -281
rect -25 -690 25 -678
<< properties >>
string FIXED_BBOX -160 -821 160 821
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2.8 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 17.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
