magic
tech sky130A
magscale 1 2
timestamp 1718126023
<< pwell >>
rect -255 -1336 255 1336
<< mvpsubdiff >>
rect -189 1258 189 1270
rect -189 1224 -81 1258
rect 81 1224 189 1258
rect -189 1212 189 1224
rect -189 1162 -131 1212
rect -189 -1162 -177 1162
rect -143 -1162 -131 1162
rect 131 1162 189 1212
rect -189 -1212 -131 -1162
rect 131 -1162 143 1162
rect 177 -1162 189 1162
rect 131 -1212 189 -1162
rect -189 -1224 189 -1212
rect -189 -1258 -81 -1224
rect 81 -1258 189 -1224
rect -189 -1270 189 -1258
<< mvpsubdiffcont >>
rect -81 1224 81 1258
rect -177 -1162 -143 1162
rect 143 -1162 177 1162
rect -81 -1258 81 -1224
<< xpolycontact >>
rect -35 684 35 1116
rect -35 -1116 35 -684
<< xpolyres >>
rect -35 -684 35 684
<< locali >>
rect -177 1224 -81 1258
rect 81 1224 177 1258
rect -177 1162 -143 1224
rect 143 1162 177 1224
rect -177 -1224 -143 -1162
rect 143 -1224 177 -1162
rect -177 -1258 -81 -1224
rect 81 -1258 177 -1224
<< viali >>
rect -19 701 19 1098
rect -19 -1098 19 -701
<< metal1 >>
rect -25 1098 25 1110
rect -25 701 -19 1098
rect 19 701 25 1098
rect -25 689 25 701
rect -25 -701 25 -689
rect -25 -1098 -19 -701
rect 19 -1098 25 -701
rect -25 -1110 25 -1098
<< properties >>
string FIXED_BBOX -160 -1241 160 1241
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 7 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 41.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
