magic
tech sky130A
magscale 1 2
timestamp 1713242186
<< metal1 >>
rect 540 -770 640 -760
rect 540 -830 550 -770
rect 630 -830 640 -770
rect 540 -840 640 -830
rect 264 -1020 270 -920
rect 370 -921 540 -920
rect 370 -1020 560 -921
rect 480 -1021 560 -1020
rect 620 -1021 810 -921
rect 540 -1110 640 -1100
rect 540 -1180 550 -1110
rect 630 -1180 640 -1110
rect 540 -1190 640 -1180
rect 540 -1400 640 -1390
rect 540 -1460 550 -1400
rect 630 -1460 640 -1400
rect 540 -1470 640 -1460
rect 710 -1550 810 -1021
rect 910 -1340 916 -1240
rect 264 -1650 270 -1550
rect 370 -1650 560 -1550
rect 620 -1650 810 -1550
rect 540 -1740 640 -1730
rect 540 -1800 550 -1740
rect 630 -1800 640 -1740
rect 540 -1810 640 -1800
<< via1 >>
rect 550 -830 630 -770
rect 270 -1020 370 -920
rect 550 -1180 630 -1110
rect 550 -1460 630 -1400
rect 810 -1340 910 -1240
rect 270 -1650 370 -1550
rect 550 -1800 630 -1740
<< metal2 >>
rect 541 -770 641 -757
rect 541 -830 550 -770
rect 630 -830 641 -770
rect 220 -920 420 -870
rect 220 -1020 270 -920
rect 370 -1020 420 -920
rect 220 -1070 420 -1020
rect 541 -1110 641 -830
rect 541 -1180 550 -1110
rect 630 -1180 641 -1110
rect 220 -1240 420 -1190
rect 541 -1240 641 -1180
rect 220 -1340 641 -1240
rect 220 -1390 420 -1340
rect 541 -1400 641 -1340
rect 760 -1240 960 -1190
rect 760 -1340 810 -1240
rect 910 -1340 960 -1240
rect 760 -1390 960 -1340
rect 541 -1460 550 -1400
rect 630 -1460 641 -1400
rect 220 -1550 420 -1500
rect 220 -1650 270 -1550
rect 370 -1650 420 -1550
rect 220 -1700 420 -1650
rect 541 -1730 641 -1460
rect 540 -1740 641 -1730
rect 540 -1800 550 -1740
rect 630 -1800 641 -1740
rect 540 -1805 641 -1800
rect 540 -1810 640 -1805
use sky130_fd_pr__nfet_01v8_648S5X  XM18
timestamp 1713229799
transform 1 0 591 0 1 -1600
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM27
timestamp 1713242186
transform 1 0 591 0 1 -971
box -211 -319 211 319
<< labels >>
flabel metal2 760 -1390 960 -1190 0 FreeSans 256 0 0 0 LO_B
port 1 nsew
flabel metal2 220 -1390 420 -1190 0 FreeSans 256 0 0 0 LO
port 3 nsew
flabel metal2 220 -1700 420 -1500 0 FreeSans 256 0 0 0 DVSS
port 6 nsew
flabel metal2 220 -1070 420 -870 0 FreeSans 256 0 0 0 DVDD
port 2 nsew
<< end >>
